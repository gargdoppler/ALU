`timescale 1 ns/1 ps
    `include "mul.v"


    module alu_tb ();
        reg clock;
        reg [31:0] a, b;
        reg [2:0] op;
        reg [31:0] correct;

        wire [31:0] out;
        wire [49:0] pro;

        alu U1 (
                .clk(clock),
                .A(a),
                .B(b),
                .OpCode(op),
                .O(out)
            );
        /* create a 10Mhz clock */
        always
        #100 clock = ~clock; // every 100 nanoseconds invert
        initial begin
            $dumpfile("alu_tb.vcd");
            $dumpvars(0,clock, a, b, op, out);
            clock = 0;

    op = 3'b011;

		/* Display the operation */
		$display ("Opcode: 011, Operation: MUL");
		/* Test Cases!*/
		a = 32'b01111000100111110001110101100111;
		b = 32'b10111000011111111111100100001001;
		correct = 32'b11110001100111110001100100010011;
		#400 //2.581786e+34 * -6.102867e-05 = -1.5756297e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110101000010001011010111010;
		b = 32'b10110101100000100000101101110001;
		correct = 32'b10110100101000111010100101111011;
		#400 //0.31462651 * -9.689085e-07 = -3.048443e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000001000111101101100100010;
		b = 32'b00111010110100001000111111111111;
		correct = 32'b10101011100001010111111000110110;
		#400 //-5.961046e-10 * 0.0015912055 = -9.485249e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110100000110101001011010000111;
		b = 32'b10010111010010100001101000000011;
		correct = 32'b01001011111101000001010011110111;
		#400 //-4.899089e+31 * -6.530255e-25 = 31992302.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011111101111000111110111000000;
		b = 32'b11100001100011110000001101100111;
		correct = 32'b11000001110100101001100101111111;
		#400 //7.982913e-20 * -3.297662e+20 = -26.32495
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011011111100010001001011110111;
		b = 32'b01110111011010110011010100101110;
		correct = 32'b11010011110111010111111001111101;
		#400 //-3.9882361e-22 * 4.7705796e+33 = -1902619800000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011111011000000111011111001100;
		b = 32'b11000001110111011110110100011010;
		correct = 32'b01100001110000101001011101010001;
		#400 //-1.6174621e+19 * -27.740772 = 4.4869648e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111010100011010100111110110111;
		b = 32'b10111101101000000100100001101011;
		correct = 32'b10111000101100001111001110011000;
		#400 //0.0010781203 * -0.07826313 = -8.437707e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101001111001000100101001011101;
		b = 32'b10111110111010101100001100100011;
		correct = 32'b10101001010100010101100111111101;
		#400 //1.0138134e-13 * -0.45852003 = -4.6485375e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011101111001101101010001010001;
		b = 32'b10110001010010010001100100110010;
		correct = 32'b11001111101101010101001101101011;
		#400 //2.079126e+18 * -2.9263671e-09 = -6084286000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000001110101011111100000011010;
		b = 32'b01011010110101110110110110001010;
		correct = 32'b01011101001101000000111011101100;
		#400 //26.746143 * 3.031878e+16 = 8.1091044e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000100010101010110010100100100;
		b = 32'b11101010101111010000001101100100;
		correct = 32'b01101111100111011000111001111111;
		#400 //-853.5803 * -1.142515e+26 = 9.752283e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010111101110100101100101111110;
		b = 32'b10100000001011001111110001010000;
		correct = 32'b10111000011110111101011110010110;
		#400 //409787060000000.0 * -1.465245e-19 = -6.0043843e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001101100110000011001010100110;
		b = 32'b10111110001111000110111110110001;
		correct = 32'b01001100011000000000111100110010;
		#400 //-319182000.0 * -0.18401982 = 58735816.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100001011001011110111000100000;
		b = 32'b10100000110110000111000101010010;
		correct = 32'b01000010110000100110011010110011;
		#400 //-2.6509144e+20 * -3.6666812e-19 = 97.200584
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011001101111101110101011001110;
		b = 32'b01010011010010100001011011010000;
		correct = 32'b01101101100101101011011001001010;
		#400 //6717302000000000.0 * 867966100000.0 = 5.8303907e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111101110111101110000011010010;
		b = 32'b11101111110110101000100010110110;
		correct = 32'b01101110001111100100001001111001;
		#400 //-0.10882725 * -1.3526601e+29 = 1.4720628e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001001011001010110111100110110;
		b = 32'b01000010111011001011010001101101;
		correct = 32'b10001100110101000010010000111010;
		#400 //-2.7617163e-33 * 118.352394 = -3.2685575e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110100000000010100011001001;
		b = 32'b00010101111111011111101000000000;
		correct = 32'b10001100111111100100101011101101;
		#400 //-3.8194453e-06 * 1.02580317e-25 = -3.917999e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011010101100010010110000000101;
		b = 32'b10110010000000101101101110110001;
		correct = 32'b10001101001101010010000011001011;
		#400 //7.32766e-23 * -7.616948e-09 = -5.5814404e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100101001110111110100100001001;
		b = 32'b01111100101101110010110110111000;
		correct = 32'b01100010100001100111010100100100;
		#400 //1.629862e-16 * 7.608941e+36 = 1.2401523e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111100011011100011011000100000;
		b = 32'b00110111001000100110101110000001;
		correct = 32'b11110100000101110010001001001001;
		#400 //-4.9474578e+36 * 9.680983e-06 = -4.7896253e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010110110011010100101001010;
		b = 32'b01010101111111000111101110100010;
		correct = 32'b11010001010101101010101111000011;
		#400 //-0.0016606238 * 34700991000000.0 = -57625293000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011110000111111101100010000011;
		b = 32'b00101100100000010000000110111011;
		correct = 32'b11001011001000010001101001011101;
		#400 //-2.879525e+18 * 3.6665926e-12 = -10558045.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101101000000110001110101011001;
		b = 32'b10001110001110000100011101011000;
		correct = 32'b10111011101111001100001101000100;
		#400 //2.536126e+27 * -2.2714102e-30 = -0.005760582
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110100001101010000001001111100;
		b = 32'b11001010011110000011100010000001;
		correct = 32'b01111111001011111000001001011100;
		#400 //-5.7364265e+31 * -4066848.2 = 2.3329176e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000111001010001000000011001001;
		b = 32'b11011101011111011110011010110110;
		correct = 32'b01100101001001110001111100100010;
		#400 //-43136.785 * -1.1434694e+18 = 4.9325594e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000111100011010101010010001111;
		b = 32'b01101100111011010011101111000110;
		correct = 32'b10110101000000101111100001001000;
		#400 //-2.126502e-34 * 2.2943815e+27 = -4.879007e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001010010011010001010111111011;
		b = 32'b11010011000111110001111000001111;
		correct = 32'b11011101111111101111000101110111;
		#400 //3360126.8 * -683404100000.0 = -2.2963244e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111110111110010000000000100100;
		b = 32'b00110000001100001010010111111000;
		correct = 32'b10101111101010111101000110000111;
		#400 //-0.4863292 * 6.4264283e-10 = -3.1253597e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000100011001111100101010100001;
		b = 32'b01001111110010001110111111000101;
		correct = 32'b10010100101101011110111101100110;
		#400 //-2.7246962e-36 * 6742313500.0 = -1.8370755e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101001000110110110110011000011;
		b = 32'b11001011110010000001100001000110;
		correct = 32'b11110101011100101111011101101010;
		#400 //1.174357e+25 * -26226828.0 = -3.0799658e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011111111100001010111011011111;
		b = 32'b00101100000010000011110011001000;
		correct = 32'b11001100100000000001011000001011;
		#400 //-3.4686089e+19 * 1.9360503e-12 = -67154010.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100111010110011101100111101;
		b = 32'b10001111011000100011000111010010;
		correct = 32'b10010100110011111101100000010011;
		#400 //1881.8512 * -1.1152255e-29 = -2.0986885e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011111100000000110111100010100;
		b = 32'b00101111011111100000010010010111;
		correct = 32'b00001111011111101110000100000111;
		#400 //5.439387e-20 * 2.3102796e-10 = 1.25665056e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011010000011001111111111001;
		b = 32'b01110001110101010000001011010001;
		correct = 32'b11111101101000010001110000111100;
		#400 //-12689401.0 * 2.1095588e+30 = -2.6769039e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011010011111000110010010111000;
		b = 32'b10110111000111100111011000001101;
		correct = 32'b00010010000111000011101010001101;
		#400 //-5.219374e-23 * -9.44502e-06 = 4.929709e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001000101011010000111010111100;
		b = 32'b00111111000000100110000110001000;
		correct = 32'b11001000001100000100011011010100;
		#400 //-354421.88 * 0.5093007 = -180507.31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011000010000011001011011000101;
		b = 32'b00110100101001110101110000000110;
		correct = 32'b11001101011111010001110111100010;
		#400 //-851413200000000.0 * 3.117313e-07 = -265412130.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101101011110101101111111010100;
		b = 32'b01110111101100110011101000011010;
		correct = 32'b01100101101011111010001101110001;
		#400 //1.42605545e-11 * 7.270309e+33 = 1.0367864e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001100001010110111100111010011;
		b = 32'b00111100001010011111110000011010;
		correct = 32'b01001000111000111011100010010011;
		#400 //44951372.0 * 0.010375047 = 466372.6
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111011110100000011110000010;
		b = 32'b10011011100101010110110100110011;
		correct = 32'b00010011100100011111000100000110;
		#400 //-1.4902909e-05 * -2.472055e-22 = 3.6840813e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011010001110111110101011100011;
		b = 32'b11101100100010000000100100010010;
		correct = 32'b01000111010001111011011011100010;
		#400 //-3.8860434e-23 * -1.315654e+27 = 51126.883
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111111110111011000111010001000;
		b = 32'b01011111000111010010001010101110;
		correct = 32'b11111111110111011000111010001000;
		#400 //nan * 1.1322804e+19 = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001110111100101100001100111001;
		b = 32'b01111111111100100000011100101111;
		correct = 32'b01111111111100100000011100101111;
		#400 //-5.98456e-30 * nan = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110011010000001000001100010110;
		b = 32'b10100010100101000000111110101100;
		correct = 32'b10010110010111101010111100100011;
		#400 //4.4822706e-08 * -4.0132074e-18 = -1.798828e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001001000000101000010110101110;
		b = 32'b00110110111011010100111010100100;
		correct = 32'b11000000011100011111101110110101;
		#400 //-534618.9 * 7.0723054e-06 = -3.780988
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011110010010110100000110000011;
		b = 32'b11000010100011011001100001001011;
		correct = 32'b00100001011000001101011111111111;
		#400 //-1.0760278e-20 * -70.79745 = 7.618002e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011101011010110000000011110010;
		b = 32'b01001110110001011101111011010110;
		correct = 32'b11101100101101011010010001001001;
		#400 //-1.05836254e+18 * 1659857700.0 = -1.7567311e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110000001101000000100010001111;
		b = 32'b10000110100111110000011110000110;
		correct = 32'b10110111010111111010110100110111;
		#400 //2.228706e+29 * -5.982021e-35 = -1.33321655e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110100010010110010000010000100;
		b = 32'b01010011011100000100111111011110;
		correct = 32'b11001000001111101010110111011011;
		#400 //-1.8917677e-07 * 1032132100000.0 = -195255.42
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110110111000101000111001101011;
		b = 32'b11011001001100101111010010010100;
		correct = 32'b11010000100111100101111101111001;
		#400 //6.7519045e-06 * -3148216400000000.0 = -21256456000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100010111001111010011100001101;
		b = 32'b01000000110001111100000100110110;
		correct = 32'b10100100001101001100000110110001;
		#400 //-6.2789547e-18 * 6.2423353 = -3.919534e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100001011001011001110011000011;
		b = 32'b00101011001001000100000110111011;
		correct = 32'b00001101000100110101001101100001;
		#400 //7.779569e-19 * 5.8355724e-13 = 4.5398236e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011011111111101110100111001110;
		b = 32'b01011110001010010000000011100011;
		correct = 32'b01111010101010000100100100111011;
		#400 //1.4350343e+17 * 3.0444957e+18 = 4.368956e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110011001100001100000111010000;
		b = 32'b00110001010011011110101000011100;
		correct = 32'b00100101000011100010110011011000;
		#400 //4.1154465e-08 * 2.9964502e-09 = 1.233173e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011110101001111100101110111001;
		b = 32'b10001111011000000010111010111000;
		correct = 32'b00101110100100101111000011100001;
		#400 //-6.0454805e+18 * -1.10530504e-29 = 6.6821e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011001010000000111000000001111;
		b = 32'b10110010100110010010100001110011;
		correct = 32'b10001100011001100100001011000010;
		#400 //9.9487974e-24 * -1.7829938e-08 = -1.7738645e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111111001111110010101111100010;
		b = 32'b11101111011100100111111110100100;
		correct = 32'b11101111001101010001011011001101;
		#400 //0.74676335 * -7.504968e+28 = -5.604435e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111001001000110110100101010111;
		b = 32'b10001011001110100011011110011000;
		correct = 32'b11000100111011011011110000001100;
		#400 //5.303006e+34 * -3.586412e-32 = -1901.8765
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010110001000001111101110001100;
		b = 32'b00010001011110011101000000011001;
		correct = 32'b10101000000111010001011110000111;
		#400 //-44250560000000.0 * 1.9706762e-28 = -8.720352e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111110001110111100111111100000;
		b = 32'b10111100011010110110001010100110;
		correct = 32'b01111011001011001011000000110010;
		#400 //-6.2411246e+37 * -0.014366781 = 8.966487e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101100010000110010000110001111;
		b = 32'b10111001001111011010010000010011;
		correct = 32'b10100110000100001000110011010111;
		#400 //2.7729795e-12 * -0.00018085567 = -5.015091e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010001010110010111100000100010;
		b = 32'b01101011010111111100010101110001;
		correct = 32'b10111101001111100001011101011111;
		#400 //-1.71553e-28 * 2.7052285e+26 = -0.046409007
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110101000000010011101100111100;
		b = 32'b11110110001000110100111011010101;
		correct = 32'b01101011101001001110000100000110;
		#400 //-4.814244e-07 * -8.280696e+32 = 3.9865296e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110001000011010110010010011011;
		b = 32'b00000100011011011101110000101000;
		correct = 32'b00110110000000110101111110111100;
		#400 //7.001442e+29 * 2.7960307e-36 = 1.9576246e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000110000100101100100100100100;
		b = 32'b01010101100111101111001000001001;
		correct = 32'b10011100001101100100010111010111;
		#400 //-2.7607323e-35 * 21845296000000.0 = -6.0309014e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000110000011100110011010000101;
		b = 32'b00100111001101001111010001101011;
		correct = 32'b00101101110010010101000000010101;
		#400 //9113.63 * 2.5112517e-15 = 2.2886618e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100101101000011101011100111011;
		b = 32'b01001100000000011001100000001110;
		correct = 32'b10110010001000111101101100101011;
		#400 //-2.8074894e-16 * 33972280.0 = -9.537682e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110001001001000101100000001000;
		b = 32'b10111101000100101001000001011011;
		correct = 32'b01101110101111000010110111000001;
		#400 //-8.1379144e+29 * -0.0357822 = 2.9119247e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110111110010000111111010101110;
		b = 32'b01000001110010101100010100011111;
		correct = 32'b00111010000111101100111001010111;
		#400 //2.3900848e-05 * 25.34625 = 0.0006057969
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001111110111111100001010001111;
		b = 32'b10011110111101100001111000100101;
		correct = 32'b10101111010101110001111101001111;
		#400 //7508139500.0 * -2.605873e-20 = -1.9565259e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011101001001101100000111110001;
		b = 32'b01001011000010111010100100010101;
		correct = 32'b00101000101101011111001011100011;
		#400 //2.2070182e-21 * 9152789.0 = 2.0200372e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000101010101001000001010010000;
		b = 32'b11001001100001001110110000111111;
		correct = 32'b01001111010111001010111011011110;
		#400 //-3400.1602 * -1088903.9 = 3702447600.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000101110110000010111110110;
		b = 32'b11011110111110001001100001101010;
		correct = 32'b01010000001101011001110100011111;
		#400 //-1.3607735e-09 * -8.956592e+18 = 12187893000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111011100000101010000101001001;
		b = 32'b10110110000100000100010101101000;
		correct = 32'b01110010000100110011110001000111;
		#400 //-1.3565397e+36 * -2.1498072e-06 = 2.9162987e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011100001000100101001010011100;
		b = 32'b01001100001010001101101100000101;
		correct = 32'b10101000110101100010001000101100;
		#400 //-5.3708074e-22 * 44264468.0 = -2.3773592e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001100110010100010111101101110;
		b = 32'b11010000110100110100100000110000;
		correct = 32'b00011110001001101101111000011011;
		#400 //-3.1151574e-31 * -28357788000.0 = 8.833897e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100111010001010110111000011001;
		b = 32'b00101000100011001011010000100110;
		correct = 32'b01010000010110010000011001001001;
		#400 //9.3233714e+23 * 1.562125e-14 = 14564271000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000110101100110011110100000111;
		b = 32'b00001000000011101110010011111000;
		correct = 32'b10001111010010000001100001010100;
		#400 //-22942.514 * 4.300072e-34 = -9.865447e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011101010011101000000111101000;
		b = 32'b10101101010110011000100011111100;
		correct = 32'b01001011001011110111101010011110;
		#400 //-9.3002686e+17 * -1.23654385e-11 = 11500190.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011000001111001001111101101101;
		b = 32'b11010010101101011000010110110010;
		correct = 32'b10101011100001011011111100111010;
		#400 //2.437892e-24 * -389816060000.0 = -9.503294e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000000100011110011101110010000;
		b = 32'b11000010110000101011011001001100;
		correct = 32'b00000011110110011110001001000100;
		#400 //-1.3153843e-38 * -97.35605 = 1.2806062e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011101011100011110010000001001;
		b = 32'b00010111011001001000011100001110;
		correct = 32'b10110101010101111110111010110100;
		#400 //-1.08937915e+18 * 7.3841236e-25 = -8.04411e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101100110001010001010101000111;
		b = 32'b11000110100111100000010001001100;
		correct = 32'b10110011111100110100110011100001;
		#400 //5.601439e-12 * -20226.148 = -1.13295535e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001010001011000110100101111010;
		b = 32'b01100101000111001010011001011101;
		correct = 32'b01101111110100110000000010100011;
		#400 //2824798.5 * 4.6234877e+22 = 1.3060421e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001111000101011010100100111111;
		b = 32'b11100010011101101101001011111001;
		correct = 32'b10110010000100000100101111111001;
		#400 //7.378863e-30 * -1.1382753e+21 = -8.399177e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100000110101110110000111000000;
		b = 32'b11000110001011111010000111100001;
		correct = 32'b10100111100100111100010000000100;
		#400 //3.6487102e-19 * -11240.47 = -4.1013217e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100001101000000001101111110111;
		b = 32'b01010011101110011110001011101110;
		correct = 32'b01110101111010001000010001000110;
		#400 //3.6918677e+20 * 1596752400000.0 = 5.8949985e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100100000101101110010011101100;
		b = 32'b01101111010000110111011110001011;
		correct = 32'b01010011111001100110110110101100;
		#400 //3.271997e-17 * 6.0494095e+28 = 1979364900000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001000100010101000110010101111;
		b = 32'b10010101010110011000001000100111;
		correct = 32'b10011110011010110110111101100010;
		#400 //283749.47 * -4.3925473e-26 = -1.246383e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011110010110011011101111101000;
		b = 32'b10111011111001011001100101011111;
		correct = 32'b11011010110000110100011110001001;
		#400 //3.9223472e+18 * -0.0070068086 = -2.7483137e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010111111001110011000100001100;
		b = 32'b11100101010001010010011010111011;
		correct = 32'b00111101101100100000101110111000;
		#400 //-1.4940406e-24 * -5.818879e+22 = 0.086936414
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000111110111001011011000001101;
		b = 32'b10010101011100001010111001010100;
		correct = 32'b00011101110011111000000011111000;
		#400 //-113004.1 * -4.8605135e-26 = 5.4925794e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101110110111110111000101011101;
		b = 32'b01000100111001010100011100000101;
		correct = 32'b01110100010010000001111001100101;
		#400 //3.4576102e+28 * 1834.2194 = 6.3420157e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110101100100100111111001011110;
		b = 32'b00101000000110001001000010110110;
		correct = 32'b10011110001011101001101110101110;
		#400 //-1.0914625e-06 * 8.469074e-15 = -9.243677e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000000010000100101111101001000;
		b = 32'b00100010101111001001100110111001;
		correct = 32'b10100011100011110011001010110000;
		#400 //-3.0370655 * 5.1120262e-18 = -1.5525558e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100000110111110001000110100001;
		b = 32'b10101001101111001100010110011111;
		correct = 32'b01001011001001000111110100100101;
		#400 //-1.28590445e+20 * -8.383159e-14 = 10779941.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111001011011011101011011110100;
		b = 32'b00101011100011110011011010100111;
		correct = 32'b01100101100001010000110111011001;
		#400 //7.7183383e+34 * 1.017593e-12 = 7.854127e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011101111011010010111111110010;
		b = 32'b10011111101100011100101100111010;
		correct = 32'b10111110001001001011101001110001;
		#400 //2.1363931e+18 * -7.5298626e-20 = -0.16086747
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000100011111011010000110111;
		b = 32'b00011000010001010100110010001010;
		correct = 32'b10001001010111011000000101001011;
		#400 //-1.045584e-09 * 2.5500296e-24 = -2.66627e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011011011000100100100010000000;
		b = 32'b00110011011101010110100010011000;
		correct = 32'b10001111010110001110101111010110;
		#400 //-1.8717708e-22 * 5.7138635e-08 = -1.06950426e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110111001001011011000000000011;
		b = 32'b00110101000111100111010000010011;
		correct = 32'b00101100110011010001101110000100;
		#400 //9.875747e-06 * 5.9028497e-07 = 5.8295053e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111000010111111101011010110010;
		b = 32'b11000011111000111011111010011001;
		correct = 32'b10111100110001110010001000000111;
		#400 //5.3367294e-05 * -455.48904 = -0.024308218
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001000001110011011001001110011;
		b = 32'b01101011000111000000110100111111;
		correct = 32'b11110011111000100110010010110100;
		#400 //-190153.8 * 1.8865498e+26 = -3.5873462e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100001010110110010111011011000;
		b = 32'b01011010010101010110001000101010;
		correct = 32'b10111100001101101011001000000110;
		#400 //-7.4262083e-19 * 1.5015526e+16 = -0.0111508425
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001001100110110010011110101101;
		b = 32'b11110101101010000000001010101110;
		correct = 32'b00111111110010111010011101010011;
		#400 //-3.7352204e-33 * -4.2595714e+32 = 1.5910438
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101011110101010000111011100110;
		b = 32'b10111001110011100100111111100101;
		correct = 32'b11100110001010111011010001111011;
		#400 //5.151431e+26 * -0.00039350908 = -2.0271349e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001110110101000000101101101000;
		b = 32'b01010100001110100000011010111110;
		correct = 32'b11100011100110100001010111011111;
		#400 //-1778758700.0 * 3195908000000.0 = -5.684749e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001100101000100111101011100110;
		b = 32'b01000001101110110100011000011110;
		correct = 32'b00001110111011011011100010001101;
		#400 //2.503402e-31 * 23.409237 = 5.8602727e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100001111000011010011111001111;
		b = 32'b01011100101110100011000100010001;
		correct = 32'b01111111001001000001111100101101;
		#400 //5.2032616e+20 * 4.1926636e+17 = 2.1815527e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111011000111110100101010001000;
		b = 32'b00001100101110011110110100110001;
		correct = 32'b10001000011001110110000011100110;
		#400 //-0.0024305899 * 2.8646518e-31 = -6.9627937e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001010001111111010011000011100;
		b = 32'b01010010001011001110001001101010;
		correct = 32'b10011101000000010110110100011011;
		#400 //-9.227557e-33 * 185633240000.0 = -1.7129414e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010110111110011100100100001101;
		b = 32'b01100101111111110110101111110110;
		correct = 32'b00111101011110010011100010011011;
		#400 //4.0355e-25 * 1.5077437e+23 = 0.060845
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101000000100110011000000010110;
		b = 32'b00010110110000010111101110111101;
		correct = 32'b10111111010111100111110011001011;
		#400 //-2.7802996e+24 * 3.1258922e-25 = -0.8690917
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110110011011101010101000001011;
		b = 32'b00000001001101000010010011101011;
		correct = 32'b00111000001001111111000111111011;
		#400 //1.2101714e+33 * 3.3087266e-38 = 4.0041265e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000001101100101000000011111101;
		b = 32'b11011110100110100110100000110000;
		correct = 32'b11100000110101110101010001111100;
		#400 //22.312983 * -5.563098e+18 = -1.241293e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000010101010101010001011111011;
		b = 32'b01011101011111000011000111110100;
		correct = 32'b01100000101010000001100110111011;
		#400 //85.31832 * 1.1357859e+18 = 9.690335e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010010011010001011111000101001;
		b = 32'b01001010001010110110111101111000;
		correct = 32'b11011101000110111101110001011101;
		#400 //-249905700000.0 * 2808798.0 = -7.019346e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101101110010110101101100010110;
		b = 32'b01001000101101111011110100000101;
		correct = 32'b11110111000100011111010001000011;
		#400 //-7.8669466e+27 * 376296.16 = -2.9603018e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111100111110000110101110001100;
		b = 32'b10110011000110011110111011011101;
		correct = 32'b01110000100101010110000000010001;
		#400 //-1.03189674e+37 * -3.5840333e-08 = 3.6983523e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100101001001101101101010011100;
		b = 32'b10011100000001011101001110101111;
		correct = 32'b01000001101011100111001100010111;
		#400 //-4.924659e+22 * -4.4279603e-22 = 21.806196
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100101101011111101011011001100;
		b = 32'b11101010001110101101011000011000;
		correct = 32'b01010000100000000101010100011110;
		#400 //-3.0503213e-16 * -5.646781e+25 = 17224495000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010100011011100100110001111110;
		b = 32'b01011001011011110100110010100110;
		correct = 32'b01101110010111101100000011000011;
		#400 //4093942200000.0 * 4209799700000000.0 = 1.7234677e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001000011110011000011101100111;
		b = 32'b01011100101110111111111110100100;
		correct = 32'b11100101101101110011111100010110;
		#400 //-255517.61 * 4.233352e+17 = -1.081696e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011101101110010000100001101001;
		b = 32'b00110011101110101001111100001000;
		correct = 32'b11010010000001101110001100001110;
		#400 //-1.6666278e+18 * 8.6902276e-08 = -144833740000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001000001111011111110100110111;
		b = 32'b10101100111011001010000110000011;
		correct = 32'b10110101101011111001110101001100;
		#400 //194548.86 * -6.725455e-12 = -1.3084295e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111111001101100000110100101100;
		b = 32'b01111111001110001101000100010001;
		correct = 32'b01111111000000110110111000100100;
		#400 //0.7111385 * 2.4566349e+38 = 1.7470075e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110100111101111101101011101000;
		b = 32'b00101000111010001111001100010010;
		correct = 32'b00011110011000011000100110111000;
		#400 //4.616661e-07 * 2.5862589e-14 = 1.193988e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011000111101011100001110001000;
		b = 32'b11110001000000100011011011111010;
		correct = 32'b11001010011110100000010000100101;
		#400 //6.352845e-24 * -6.447922e+29 = -4096265.2
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001001000100110100001100111010;
		b = 32'b10000010111001010000101001111110;
		correct = 32'b00001100100000111100000100101100;
		#400 //-603187.6 * -3.3654548e-37 = 2.0300007e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110001101100000111001101111100;
		b = 32'b10100101100100110010101100100111;
		correct = 32'b00010111110010101110000000011101;
		#400 //-5.135403e-09 * -2.5529676e-16 = 1.3110518e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100001010100110101001011000100;
		b = 32'b11111000010001100110011101111011;
		correct = 32'b01011010001000111100011101101111;
		#400 //-7.159912e-19 * -1.6096463e+34 = 1.1524925e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010000111010010011010001011001;
		b = 32'b00001000011001011001111011001100;
		correct = 32'b00011001110100010010110001111100;
		#400 //31300176000.0 * 6.9098846e-34 = 2.162806e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100001001100101011000011110111;
		b = 32'b01001111100111101001110100011010;
		correct = 32'b10110001010111010110110111000010;
		#400 //-6.0542957e-19 * 5322192000.0 = -3.2222123e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011000000111101010110010110110;
		b = 32'b11011011100011101101000010101000;
		correct = 32'b01110100001100010000101001000011;
		#400 //-697858500000000.0 * -8.039773e+16 = 5.6106242e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011000100001101111011100011110;
		b = 32'b11101111101011110010011011011100;
		correct = 32'b01001000101110001010111011010100;
		#400 //-3.4887713e-24 * -1.0841371e+29 = 378230.62
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000001001001011100100001000011;
		b = 32'b00100001000010010001011001001010;
		correct = 32'b10100010101100011000110100110110;
		#400 //-10.361392 * 4.6446905e-19 = -4.812546e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000111101111001001101100101110;
		b = 32'b00111110101100100010101111001100;
		correct = 32'b10000111000000110100010000101010;
		#400 //-2.8378302e-34 * 0.3479904 = -9.875376e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011110000000011011011111011100;
		b = 32'b11000101101100001001010011011000;
		correct = 32'b11100100001100101111001110100110;
		#400 //2.3367954e+18 * -5650.6055 = -1.3204309e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011100101100001101111000111111;
		b = 32'b01111000010101001111000001111110;
		correct = 32'b01010101100100110001111000110100;
		#400 //1.1704152e-21 * 1.7275698e+34 = 20219741000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001110010111110111100011111001;
		b = 32'b10111101010111111001111110110011;
		correct = 32'b00001100010000110011010111001001;
		#400 //-2.7545118e-30 * -0.05459566 = 1.5038439e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010010111111001011100110110110;
		b = 32'b10000111011010001111010110100111;
		correct = 32'b10011010111001011111101011010000;
		#400 //542723740000.0 * -1.7525931e-34 = -9.511739e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010100110100011010011010101101;
		b = 32'b01111010110110111011000111010101;
		correct = 32'b01010000001100111110101100111001;
		#400 //2.1169349e-26 * 5.7035994e+35 = 12074149000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100000010011000001101011100010;
		b = 32'b00001101010110101001111010010010;
		correct = 32'b10101110001011100100110101010001;
		#400 //-5.8829264e+19 * 6.736731e-31 = -3.963169e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011111011111111100110101001011;
		b = 32'b00111100101000100000001110110111;
		correct = 32'b11011100101000011110001110100000;
		#400 //-1.8432471e+19 * 0.019777162 = -3.6454198e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110000011011010110100010110;
		b = 32'b11011100100101111111001101110110;
		correct = 32'b11011011001010000010111110101001;
		#400 //0.13835558 * -3.4216328e+17 = -4.73402e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111000000111111101110011101110;
		b = 32'b10101001001001111111110011100010;
		correct = 32'b11100001110100011100111000010100;
		#400 //1.2969628e+34 * -3.730079e-14 = -4.8377738e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101000010100010000111000001010;
		b = 32'b10110111001001010111000111110111;
		correct = 32'b11100000000001110001101100011101;
		#400 //3.9489343e+24 * -9.861301e-06 = -3.8941628e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101110110100111111001011000010;
		b = 32'b00101000100101011010000110001011;
		correct = 32'b01010111111101111100010000010011;
		#400 //3.2797407e+28 * 1.6612381e-14 = 544843000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100111001000100011111000001101;
		b = 32'b00111111100111111100101100100110;
		correct = 32'b01100111010010101000101010010011;
		#400 //7.66168e+23 * 1.2483871 = 9.564743e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110110000101110101011110011110;
		b = 32'b01000110010011110000111000111011;
		correct = 32'b00111100111101001101000010000101;
		#400 //2.2551753e-06 * 13251.558 = 0.029884586
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001111110110100110001100111111;
		b = 32'b11001001000011101011011000111110;
		correct = 32'b01011001011100110111110100001001;
		#400 //-7327874600.0 * -584547.9 = 4283493600000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100001011101001111101101110101;
		b = 32'b11101001000011101001000101011001;
		correct = 32'b11001011000010000110111010010010;
		#400 //8.3003216e-19 * -1.0772116e+25 = -8941202.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011100100101100101011100001100;
		b = 32'b11011010011100001001110101101111;
		correct = 32'b10110111100011010100111000010000;
		#400 //9.948668e-22 * -1.6931774e+16 = -1.684486e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111110000010111100101001011010;
		b = 32'b00100011010011100101100010010001;
		correct = 32'b01100001111000010101101001100010;
		#400 //4.645334e+37 * 1.1186037e-17 = 5.1962877e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101000110101101010000110101010;
		b = 32'b10011110010010100001011011110110;
		correct = 32'b11000111101010010110111011010000;
		#400 //8.108549e+24 * -1.0698539e-20 = -86749.625
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010011010111100001010001110101;
		b = 32'b00011101111110011110100011011001;
		correct = 32'b10110001110110001100101111100101;
		#400 //-953825950000.0 * 6.615051e-21 = -6.3096075e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001010100010001100010111111100;
		b = 32'b11010111110001001100100000001010;
		correct = 32'b10100010110100100100010011101010;
		#400 //1.3170797e-32 * -432726880000000.0 = -5.699358e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010111011101011100001011110111;
		b = 32'b11011111101011111100111100100110;
		correct = 32'b00110111101010001100011100100100;
		#400 //-7.940985e-25 * -2.5336772e+19 = 2.0119893e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101001110101111110100000110101;
		b = 32'b10000010000001110001001101001000;
		correct = 32'b00101100011000111101011101101110;
		#400 //-3.2626952e+25 * -9.923767e-38 = 3.2378228e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101011100110000111100111110010;
		b = 32'b11000111000111101001101011110010;
		correct = 32'b11110011001111001110111100011010;
		#400 //3.686652e+26 * -40602.945 = -1.4968893e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100111101000010001001011011010;
		b = 32'b00011011101101000000111111100000;
		correct = 32'b11000011111000101001011001111101;
		#400 //-1.5212975e+24 * 2.978876e-22 = -453.1757
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010000001011100110110111001100;
		b = 32'b01001011110100000100010001111001;
		correct = 32'b00011100100011011110011111011101;
		#400 //3.4400034e-29 * 27298034.0 = 9.390533e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010010110111000101000011010110;
		b = 32'b01010001100101101111100000101010;
		correct = 32'b10100101000000011110110011110000;
		#400 //-1.390388e-27 * 81051075000.0 = -1.1269244e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000111010100001110101010100111;
		b = 32'b11110011110100001001111000110010;
		correct = 32'b10111011101010100011111111000001;
		#400 //1.5717139e-34 * -3.3056834e+31 = -0.0051955883
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010100101100101001011010110001;
		b = 32'b11100010011011001001000101011110;
		correct = 32'b11110111101001010000100001010100;
		#400 //6136259000000.0 * -1.0909766e+21 = -6.694515e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010000101101101001100111011100;
		b = 32'b10111111111101010011101001010111;
		correct = 32'b11010001001011101110101011011100;
		#400 //24508293000.0 * -1.9158429 = -46954037000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010111100000100110111001110000;
		b = 32'b11011110101001011110001010101101;
		correct = 32'b01110110101010010000100101011000;
		#400 //-286821670000000.0 * -5.9766533e+18 = 1.7142338e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111000001110100100011110001000;
		b = 32'b10010101101001101101001000001000;
		correct = 32'b11001110011100101100011001101101;
		#400 //1.5112782e+34 * -6.737824e-26 = -1018272600.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001111000000111001001011110011;
		b = 32'b10100100100011111011110101011011;
		correct = 32'b00110100000100111100000011010000;
		#400 //-2207445800.0 * -6.2337145e-17 = 1.3760587e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101000011100000011000001101100;
		b = 32'b11100001001111010101000101011101;
		correct = 32'b01001010001100011010000000010110;
		#400 //-1.3333176e-14 * -2.182686e+20 = 2910213.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100011101010100000000110001011;
		b = 32'b01111110110101110010010000100010;
		correct = 32'b01100011000011101101111101001011;
		#400 //1.843209e-17 * 1.4298582e+38 = 2.6355276e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000101111011000111001111100110;
		b = 32'b11000011111100101111101100111011;
		correct = 32'b10001010011000000110110110011100;
		#400 //2.2235908e-35 * -485.96274 = -1.0805823e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100001001100000000011111101100;
		b = 32'b11101000000100000100001000010110;
		correct = 32'b11001001110001100110001111001100;
		#400 //5.9641604e-19 * -2.7249594e+24 = -1625209.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110110111011101011100011110;
		b = 32'b00101011110100010101011010000010;
		correct = 32'b00101011001101010110011110010110;
		#400 //0.43328184 * 1.4874354e-12 = 6.444787e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001100011001100100010100011011;
		b = 32'b00000111110000111000101011101011;
		correct = 32'b00010100101011111110001110011000;
		#400 //60363884.0 * 2.9421988e-34 = 1.7760254e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001010110111111010110101001110;
		b = 32'b01110100111001110111100000011001;
		correct = 32'b11000000010010100011111001010000;
		#400 //-2.1539309e-32 * 1.4671099e+32 = -3.1600533
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100100011010110000000010100101;
		b = 32'b10010111001100011011111010001010;
		correct = 32'b00111100001000110010101001011011;
		#400 //-1.7340125e+22 * -5.743228e-25 = 0.009958829
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011001011011110011001010110101;
		b = 32'b01000100100110100110101110011110;
		correct = 32'b11011110100100000100100100001111;
		#400 //-4208017000000000.0 * 1235.363 = -5.198429e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011100000011010110000100000101;
		b = 32'b11100010000111011001011001001100;
		correct = 32'b01111110101011100000111100000010;
		#400 //-1.5917858e+17 * -7.267422e+20 = 1.156818e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010111111001001110100000100111;
		b = 32'b11101100001000001001011010001100;
		correct = 32'b11000100100011111001011110110110;
		#400 //1.4792758e-24 * -7.765563e+26 = -1148.741
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000011101101111111011111111000;
		b = 32'b11100010011101111010110011010100;
		correct = 32'b10100110101100011111110001110011;
		#400 //1.0812704e-36 * -1.14219984e+21 = -1.2350269e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010101001101010100101011110111;
		b = 32'b00110011010001000101010111010011;
		correct = 32'b11001001000010110000101000101100;
		#400 //-12458349000000.0 * 4.5712863e-08 = -569506.75
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101111100001110011000100101011;
		b = 32'b01010110001000010101001000001011;
		correct = 32'b01000110001010100110001001111111;
		#400 //2.4591293e-10 * 44343436000000.0 = 10904.624
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000010101110011100011010100001;
		b = 32'b01011111100010101000111011011111;
		correct = 32'b01100010110010010001100110000010;
		#400 //92.88795 * 1.9968325e+19 = 1.8548168e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011110101100111100111001101010;
		b = 32'b11110001010110000010011100001111;
		correct = 32'b11010000100101111101000110011000;
		#400 //1.9037733e-20 * -1.0703357e+30 = -20376764000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010100011101000110001011101101;
		b = 32'b11111110111000001000111100001101;
		correct = 32'b11010011110101100101111100011111;
		#400 //1.23383616e-26 * -1.4924492e+38 = -1841437700000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111011110001101001101111101010;
		b = 32'b11001110101100101111100111011111;
		correct = 32'b01001011000010101101101001000011;
		#400 //-0.006061067 * -1501360000.0 = 9099843.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101000010011110110111011001100;
		b = 32'b11010011010000010110110100000000;
		correct = 32'b11111100000111001011101011011010;
		#400 //3.9182948e+24 * -830757400000.0 = -3.2551524e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100000011001111001011100001001;
		b = 32'b00100100001111001100010010111111;
		correct = 32'b11000101001010101100010011100111;
		#400 //-6.6751267e+19 * 4.0932652e-17 = -2732.3064
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011111111001111101100011011;
		b = 32'b00001111001110100110000010001001;
		correct = 32'b10011011101110000010110111010111;
		#400 //-33158710.0 * 9.1891e-30 = -3.046987e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010101001101000010011001001100;
		b = 32'b11011110100010111010011000101100;
		correct = 32'b10110100010001001000101101110110;
		#400 //3.638092e-26 * -5.0313894e+18 = -1.8304658e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100011100011001001010110001000;
		b = 32'b11111110001100100010011110011001;
		correct = 32'b11100010010000111010101101101111;
		#400 //1.524216e-17 * -5.9202047e+37 = -9.0236705e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011110011110101110101110110000;
		b = 32'b11011100011011001110111100001010;
		correct = 32'b01111011011010000011101110010010;
		#400 //-4.5201847e+18 * -2.6676368e+17 = 1.2058211e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100010111001010100011111011110;
		b = 32'b10100001101000100000011000011000;
		correct = 32'b01000101000100010001110011110000;
		#400 //-2.1147415e+21 * -1.097916e-18 = 2321.8086
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110001110100001111111010101101;
		b = 32'b00101010110111110110010110110100;
		correct = 32'b10011101001101100110000011100000;
		#400 //-6.08255e-09 * 3.9683328e-13 = -2.4137583e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011111111000101000101010111010;
		b = 32'b00111111011110100100001100011110;
		correct = 32'b11011111110111010111011011011110;
		#400 //-3.2648129e+19 * 0.9775866 = -3.1916373e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000000001010100100000110100001;
		b = 32'b10011101001110001101100111101110;
		correct = 32'b00011101111101011110000000110111;
		#400 //-2.6602557 * -2.4464864e-21 = 6.5082793e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000100000101001111011000100001;
		b = 32'b11011010100101011010001001111001;
		correct = 32'b10011111001011100010001110010111;
		#400 //1.7510333e-36 * -2.1059206e+16 = -3.6875372e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100001100101110110001010111110;
		b = 32'b10101001111011001110000010100101;
		correct = 32'b01001100000011000001001111011111;
		#400 //-3.490717e+20 * -1.0519475e-13 = 36720508.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100010011000000011100100000;
		b = 32'b10000000110111100000110000011110;
		correct = 32'b10000101101100001111011111010110;
		#400 //816.1113 * -2.0391827e-38 = -1.6642001e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001011000010001001100011101010;
		b = 32'b11110000101001101000100101110110;
		correct = 32'b10111100001100011011100100000001;
		#400 //2.6307687e-32 * -4.1232553e+29 = -0.010847331
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100101001011100101110010011110;
		b = 32'b00110101000001111100010100110110;
		correct = 32'b01011010101110001111001001010011;
		#400 //5.1462516e+22 * 5.05784e-07 = 2.6028917e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000011001110011001000010011;
		b = 32'b00011001101001010101001010010011;
		correct = 32'b10001010100101010100110111011001;
		#400 //-8.410847e-10 * 1.7093952e-23 = -1.4377461e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010001000110101010100001110100;
		b = 32'b00100010100101110100000111110000;
		correct = 32'b10110100001101101100001001100100;
		#400 //-41515696000.0 * 4.0998446e-18 = -1.702079e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000001101000000111110100001111;
		b = 32'b00000101011100010100100100000011;
		correct = 32'b10000111100101110100001110000001;
		#400 //-20.061064 * 1.1345176e-35 = -2.275963e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001010011101111110011000101001;
		b = 32'b00101111100100100100100110000100;
		correct = 32'b10111010100011011010100001110100;
		#400 //-4061578.2 * 2.660948e-10 = -0.0010807649
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100100111001110101000010100111;
		b = 32'b11011001001111001001001010100110;
		correct = 32'b10111110101010100110001110111101;
		#400 //1.0031691e-16 * -3317408600000000.0 = -0.3327922
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110100001100010001010000001100;
		b = 32'b11001000101000001011000000100110;
		correct = 32'b10111101010111100100110010111111;
		#400 //1.6491703e-07 * -329089.2 = -0.05427241
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100001110000110010010101100010;
		b = 32'b10101101000010110111000101010101;
		correct = 32'b11001111010101001001011101100001;
		#400 //4.499761e+20 * -7.9264e-12 = -3566690600.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101001001001011011010011110001;
		b = 32'b11001000111100010101111110001100;
		correct = 32'b11110010100111000011110100110000;
		#400 //1.2520452e+25 * -494332.38 = -6.189265e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001101110011101011101111000001;
		b = 32'b01010101001111010011010011000010;
		correct = 32'b01100011100110001100101100111000;
		#400 //433551400.0 * 13002143000000.0 = 5.637097e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110001110111000000011001111000;
		b = 32'b01010001010111001011110100110000;
		correct = 32'b11000011101111011011100000101001;
		#400 //-6.403578e-09 * 59254178000.0 = -379.43875
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100000100100001100110100000011;
		b = 32'b10011111011100111001010100100110;
		correct = 32'b00000000100010011100011011110111;
		#400 //-2.4530214e-19 * -5.1580624e-20 = 1.2652838e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101101001001100110011100000011;
		b = 32'b00101011000101101101011001111011;
		correct = 32'b11011000110001000001011110001100;
		#400 //-3.2186903e+27 * 5.3588357e-13 = -1724843300000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100110010111000100111110010111;
		b = 32'b10110101110101100111100101000101;
		correct = 32'b11011100101110001001001011100101;
		#400 //2.600972e+23 * -1.5979537e-06 = -4.1562326e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011001100111111010010010010001;
		b = 32'b10001001111100100000001011100111;
		correct = 32'b00100100000101101110101101100000;
		#400 //-5616933000000000.0 * -5.826211e-33 = 3.2725436e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010000111010011000101001111100;
		b = 32'b10000110010110101101111101111000;
		correct = 32'b10010111110001111010101111001011;
		#400 //31345336000.0 * -4.1165422e-35 = -1.290344e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110100110111000010110000011100;
		b = 32'b10011000011011111001110100111010;
		correct = 32'b01001101110011100001010001100111;
		#400 //-1.3955078e+32 * -3.0969405e-24 = 432180450.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011000000100010110011100011101;
		b = 32'b01010001100101101101100110111001;
		correct = 32'b11101010001010110101110000101001;
		#400 //-639488200000000.0 * 80987234000.0 = -5.179038e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000100010000110010010010101110;
		b = 32'b11100000001011001010101010101100;
		correct = 32'b00100101000000111001111010111110;
		#400 //-2.2938982e-36 * -4.9767784e+19 = 1.1416223e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001101111001000001011001111011;
		b = 32'b11011001001011011000110001001001;
		correct = 32'b00100111100110101010000000101110;
		#400 //-1.4056997e-30 * -3053088500000000.0 = 4.2917254e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001001100110101001110010011100;
		b = 32'b11001101101000110011110110100010;
		correct = 32'b11010111110001010010110111100001;
		#400 //1266579.5 * -342340670.0 = -433601680000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100100101100000011001110001010;
		b = 32'b01110101010100000111111101110010;
		correct = 32'b01011010100011111000000110011000;
		#400 //7.6415144e-17 * 2.643024e+32 = 2.0196706e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010101010101111101101101011000;
		b = 32'b10111001100001101001010001010010;
		correct = 32'b00001111011000101111001111000000;
		#400 //-4.3591936e-26 * -0.0002566898 = 1.1189605e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001011101001101010000001001111;
		b = 32'b11010110001100100010010101111001;
		correct = 32'b10100010011001111110011110110110;
		#400 //6.418208e-32 * -48968503000000.0 = -3.1429004e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000001011110100010001011010110;
		b = 32'b10000101111011010100110000011001;
		correct = 32'b00000111111001111101110010011011;
		#400 //-15.633505 * -2.2315327e-35 = 3.4886677e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000011100000001101110111101100;
		b = 32'b10010011001011110001111000110001;
		correct = 32'b00010111001100000100110111001110;
		#400 //-257.73376 * -2.210299e-27 = 5.696687e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111011101001100010011010001000;
		b = 32'b01001100100100110010011011100111;
		correct = 32'b11001000101111110000001010111111;
		#400 //-0.0050705113 * 77150010.0 = -391189.97
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101110111101011001010000110111;
		b = 32'b10100011010101000100101011000101;
		correct = 32'b01010010110010111010011001110111;
		#400 //-3.8001504e+28 * -1.1508376e-17 = 437335600000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110000001011101100110111111001;
		b = 32'b01101010110101000101100111110111;
		correct = 32'b01011011100100010000000000000000;
		#400 //6.3593536e-10 * 1.2835856e+26 = 8.162774e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011010111100101101111101001110;
		b = 32'b01101111111111101010010111101110;
		correct = 32'b11001011011100011001011011111011;
		#400 //-1.0044962e-22 * 1.5761958e+29 = -15832827.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110110001000101111001000110010;
		b = 32'b10010100110001010000111010010101;
		correct = 32'b11001011011110101101101101010001;
		#400 //8.262348e+32 * -1.9897668e-26 = -16440145.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001101001011101011010100111101;
		b = 32'b10101001001100010000111111010111;
		correct = 32'b00110110111100011010110000111101;
		#400 //-183194580.0 * -3.9315634e-14 = 7.202411e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010110000111000010011101111010;
		b = 32'b00000100100001010101111100110100;
		correct = 32'b10011011001000101011010100101010;
		#400 //-42923340000000.0 * 3.135558e-36 = -1.3458863e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000010010011011000011111111111;
		b = 32'b10111101101000100011000010001000;
		correct = 32'b01000000100000100011011100000110;
		#400 //-51.38281 * -0.07919413 = 4.0692167
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001100000000010100110011001010;
		b = 32'b10111101101010100110010101010110;
		correct = 32'b10001010001011000010000001011010;
		#400 //9.960906e-32 * -0.083201095 = -8.2875834e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011001001111100110010110110100;
		b = 32'b01111000010101000010010110010110;
		correct = 32'b01010010000111011100100000101101;
		#400 //9.8433086e-24 * 1.7211395e+34 = 169417060000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100100000101111011101000110001;
		b = 32'b10110001001110000010010100011000;
		correct = 32'b11010101110110100100011110011111;
		#400 //1.11955e+22 * -2.679661e-09 = -30000143000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101011110010011100101111110110;
		b = 32'b10110000110000011110011011001110;
		correct = 32'b00011101000110001101100010110100;
		#400 //-1.433852e-12 * -1.4108197e-09 = 2.0229065e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111010001111000000100001010000;
		b = 32'b10111000001100001000011111001000;
		correct = 32'b01110011000000011010100101110010;
		#400 //-2.440801e+35 * -4.2088126e-05 = 1.0272874e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011110000001111101001100101010;
		b = 32'b11000001111000110101000100100100;
		correct = 32'b01100000011100010011011010010110;
		#400 //-2.4468031e+18 * -28.41462 = 6.952498e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111111100110000110101101101;
		b = 32'b01000001110000101001111011101011;
		correct = 32'b10111010001110001100011100001110;
		#400 //-2.897411e-05 * 24.327597 = -0.00070487044
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010010111111110010000000101101;
		b = 32'b01001101111001001100110100001101;
		correct = 32'b00100001011001000000010100000010;
		#400 //1.6100694e-27 * 479830430.0 = 7.725603e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000000111111000011011010010100;
		b = 32'b11001100111111001111100110100001;
		correct = 32'b11001110011110010011101110101001;
		#400 //7.8816624 * -132631816.0 = -1045359170.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001010001010101010000011001111;
		b = 32'b01111000101000000100010011011011;
		correct = 32'b11000011010101011010010011001100;
		#400 //-8.215447e-33 * 2.6005127e+34 = -213.64374
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101100010011000000101110110101;
		b = 32'b10010010001101101100010111000000;
		correct = 32'b00111111000100011010110111110001;
		#400 //-9.867046e+26 * -5.767282e-28 = 0.5690604
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111001010011111011010000010100;
		b = 32'b01111001010101111101010110010101;
		correct = 32'b01110011001011110001110110000111;
		#400 //0.00019808143 * 7.0042236e+34 = 1.3874067e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111111010111100100010010000011;
		b = 32'b10101010010111011011001111001100;
		correct = 32'b00101010010000000111110101000000;
		#400 //-0.8682329 * -1.9691123e-13 = 1.709648e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100100110101010010100000011000;
		b = 32'b01001101110110100111011011010000;
		correct = 32'b01110011001101011110011100010010;
		#400 //3.1456364e+22 * 458152450.0 = 1.441181e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011111100110011100101100000011;
		b = 32'b00111100101000010011011101110011;
		correct = 32'b11011100110000011011001111111001;
		#400 //-2.216391e+19 * 0.01967976 = -4.3618042e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100000000111001000100111000111;
		b = 32'b11001110010011101000111001111110;
		correct = 32'b10101110111111001001101111111111;
		#400 //1.3259301e-19 * -866361200.0 = -1.1487344e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101101100111001000111001010101;
		b = 32'b01001001010010011010011011011100;
		correct = 32'b11110111011101101010001110010111;
		#400 //-6.0564663e+27 * 825965.75 = -5.0024337e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111111100101111001110101111001;
		b = 32'b01111101110101000011000010100000;
		correct = 32'b01111101111110110101011001101001;
		#400 //1.1844932 * 3.5256101e+37 = 4.1760612e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101010010000111110011010011111;
		b = 32'b10111010101001111001101100011101;
		correct = 32'b00100101100000000100001000100101;
		#400 //-1.7399492e-13 * -0.0012787316 = 2.2249282e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001100001110100100001111100110;
		b = 32'b01100110100010000101110001010110;
		correct = 32'b00110011010001100110111010000010;
		#400 //1.4349351e-31 * 3.2197257e+23 = 4.6200974e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101010110010111011011110110111;
		b = 32'b11111101110100001111011111101011;
		correct = 32'b11101001001001100100101010001110;
		#400 //3.6187522e-13 * -3.4720836e+37 = -1.256461e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010011101101100011001000111001;
		b = 32'b01000101001011011110111111110011;
		correct = 32'b01011001011101111001010101101101;
		#400 //1565053300000.0 * 2782.9968 = 4355538400000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110101111100111110101101000010;
		b = 32'b11111101111011001000011001011000;
		correct = 32'b01110100011000010101110011100010;
		#400 //-1.817338e-06 * -3.929942e+37 = 7.142033e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000001001101111011000011110111;
		b = 32'b01000110100010010100111011011010;
		correct = 32'b11001000010001010000110010010001;
		#400 //-11.480704 * 17575.426 = -201778.27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101111111101101111011101000010;
		b = 32'b01101111110100101111111110010000;
		correct = 32'b11100000010010111000110101011111;
		#400 //-4.4922827e-10 * 1.3060162e+29 = -5.8669936e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110010101000010011101010010011;
		b = 32'b11101000000111000000101101101011;
		correct = 32'b01011011010001001000110111000101;
		#400 //-1.8769503e-08 * -2.9475992e+24 = 5.5324973e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001111011100110001111010100111;
		b = 32'b00100000111100000100010010110101;
		correct = 32'b10110000111001000010110111111101;
		#400 //-4078872300.0 * 4.0703048e-19 = -1.6602254e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000001110111100101000101000100;
		b = 32'b00111001100110001111011000100011;
		correct = 32'b10111100000001001101011000000001;
		#400 //-27.78968 * 0.00029175085 = -0.008107663
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100010100011111001110110100101;
		b = 32'b00000011010101101111110101101000;
		correct = 32'b00100110011100010011011111100010;
		#400 //1.324622e+21 * 6.3179844e-37 = 8.3689407e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111100001001011011011010010011;
		b = 32'b01000000110000101010110111100000;
		correct = 32'b00111101011111000000100111010010;
		#400 //0.01011433 * 6.083725 = 0.061532803
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010111110011001011101010001000;
		b = 32'b10001101000010010010100010011101;
		correct = 32'b10100101010110110110000010011011;
		#400 //450203040000000.0 * -4.226527e-31 = -1.9027953e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100101110000101001010101010101;
		b = 32'b00010111111110001001011000000110;
		correct = 32'b00111110001111001111001010110010;
		#400 //1.1486172e+23 * 1.6064496e-24 = 0.18451956
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000011000010101010000111000111;
		b = 32'b01111011110011000111001101111110;
		correct = 32'b01111111010111010110111011101011;
		#400 //138.63194 * 2.123142e+36 = 2.943353e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000011010011110010001100100011;
		b = 32'b01011110000110001001001101011100;
		correct = 32'b10100001111101101110100000110001;
		#400 //-6.0872168e-37 * 2.748558e+18 = -1.6731069e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001100011100111001100110011001;
		b = 32'b11010000000000010111011000100101;
		correct = 32'b10011100111101100110000110100100;
		#400 //1.8766261e-31 * -8688014000.0 = -1.6304154e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100000110111110011101111011101;
		b = 32'b10110101100110100111110111111110;
		correct = 32'b00010111000001101011011111100001;
		#400 //-3.7817284e-19 * -1.1510563e-06 = 4.3529823e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010100011111001010011010110110;
		b = 32'b11001110101110011100110001001000;
		correct = 32'b10100011101101110101111000010101;
		#400 //1.27556266e-26 * -1558586400.0 = -1.9880745e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000101110100000010111100110010;
		b = 32'b11011010000101101101010111100100;
		correct = 32'b00100000011101010101001100110000;
		#400 //-1.9577563e-35 * -1.0614105e+16 = 2.0779832e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000111000000010011000001101011;
		b = 32'b11111011110000111000011000010011;
		correct = 32'b01000011010001010101011100010101;
		#400 //-9.71911e-35 * -2.0304345e+36 = 197.34016
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100110101000100000110100000101;
		b = 32'b10110111011000100101111001111110;
		correct = 32'b01011110100011110100101101001111;
		#400 //-3.8263177e+23 * -1.349265e-05 = 5.1627167e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101001011000011001111000111101;
		b = 32'b10100101101101000011001111010010;
		correct = 32'b00001111100111101101000011101110;
		#400 //-5.0097286e-14 * -3.1260137e-16 = 1.566048e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100110111101111111011100010001;
		b = 32'b10110111110111011010010001010111;
		correct = 32'b10011111010101101010111101111000;
		#400 //1.7206035e-15 * -2.642178e-05 = -4.5461407e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111011011011011101001001001100;
		b = 32'b00000000111101011110110111100001;
		correct = 32'b10111100111001000111011100111111;
		#400 //-1.2348397e+36 * 2.2585031e-38 = -0.027888892
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000001101111110010000000100001;
		b = 32'b10010110100110001011011110100101;
		correct = 32'b00011000111001000000100001011101;
		#400 //-23.890688 * -2.467282e-25 = 5.8945063e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000011110000000000001010000000;
		b = 32'b11110111100101100100001111111100;
		correct = 32'b11111011111000010110100011101001;
		#400 //384.01953 * -6.0954954e+33 = -2.3407892e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100010110110001010101111000010;
		b = 32'b10011010010111000111011101001010;
		correct = 32'b00111101101110101001100010010001;
		#400 //-1.9984366e+21 * -4.5591295e-23 = 0.09111131
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000010101111001010010101011010;
		b = 32'b10110100110110111111110110011110;
		correct = 32'b00111000001000100001110001011000;
		#400 //-94.32295 * -4.097646e-07 = 3.8650207e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001110000111000011001011011001;
		b = 32'b11101000101000001100110110101100;
		correct = 32'b01110111010001000011101010001011;
		#400 //-655144500.0 * -6.074981e+24 = 3.9799905e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010110110110110001011100001000;
		b = 32'b01011010101011100010000011110100;
		correct = 32'b10110010000101010000010111011011;
		#400 //-3.5395893e-25 * 2.450644e+16 = -8.674273e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110110011110110111110110101110;
		b = 32'b00111001111000001101101100100010;
		correct = 32'b01110000110111001110010100111110;
		#400 //1.27521055e+33 * 0.00042887876 = 5.469107e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110010001101111111001010000001;
		b = 32'b00010111000110101010101101110111;
		correct = 32'b00001001110111100100011000101100;
		#400 //1.0707141e-08 * 4.9976503e-25 = 5.3510545e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101110010010001101101010100010;
		b = 32'b10010101101011100011100011011101;
		correct = 32'b10000100100010001011000100110111;
		#400 //4.566892e-11 * -7.0367755e-26 = -3.2136192e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011111100111110000101110111111;
		b = 32'b10111101100111101101110110110000;
		correct = 32'b11011101110001010110010111110101;
		#400 //2.2920927e+19 * -0.07757127 = -1.7780055e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010100111010110110010001110010;
		b = 32'b10001001001010110011001101111101;
		correct = 32'b00011110100111010110101101110000;
		#400 //-8088020000000.0 * -2.0607586e-33 = 1.6667457e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011011010001110100010010111001;
		b = 32'b11010100101000011001101110011111;
		correct = 32'b00110000011110111001011010110101;
		#400 //-1.64831e-22 * -5552805000000.0 = 9.1527436e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010100010010110110000000100001;
		b = 32'b11100111010110011010101110100001;
		correct = 32'b01111100001011001110110011010101;
		#400 //-3493964500000.0 * -1.0279195e+24 = 3.5915143e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100101110000001100110011010111;
		b = 32'b10001010010010101010111001101010;
		correct = 32'b00110000100110001010010011111101;
		#400 //-1.1380912e+23 * -9.75875e-33 = 1.1106348e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000101010111101001000010101101;
		b = 32'b00110110110011101110011110001000;
		correct = 32'b10111100101100111110000110110110;
		#400 //-3561.0422 * 6.166232e-06 = -0.021958213
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011111011101010110011110000101;
		b = 32'b11101111010010110010110010001101;
		correct = 32'b11001111010000101100001111001011;
		#400 //5.1966397e-20 * -6.2879316e+28 = -3267611400.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000111101101010111111110101011;
		b = 32'b11010110110110100111110011101000;
		correct = 32'b10011111000110101110011101000110;
		#400 //2.730889e-34 * -120115000000000.0 = -3.2802073e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010110011100101001111111001001;
		b = 32'b10111101010001100001110111110110;
		correct = 32'b00010100001110111100001111111011;
		#400 //-1.9599024e-25 * -0.048368417 = 9.479738e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111101111000000111001110010111;
		b = 32'b10001010111000001101010101011100;
		correct = 32'b10001001010001010010000000110101;
		#400 //0.10959547 * -2.1650672e-32 = -2.3728156e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010010011111100010001000011110;
		b = 32'b10111100010011010011010010001110;
		correct = 32'b00001111010010111011010101111110;
		#400 //-8.019032e-28 * -0.012524737 = 1.0043627e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011110010010111111110111111001;
		b = 32'b10010011010011000001001100101001;
		correct = 32'b10110010001000101001110110100111;
		#400 //3.6747946e+18 * -2.5757867e-27 = -9.465487e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100011100101110101110000101100;
		b = 32'b00110011110001000100001110010101;
		correct = 32'b00010111111010000001010100001110;
		#400 //1.6410489e-17 * 9.139254e-08 = 1.4997964e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101001101010011111100110111111;
		b = 32'b01101001011110000001011110000010;
		correct = 32'b01010011101001001011100110001101;
		#400 //7.548432e-14 * 1.8745288e+25 = 1414975300000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110011000001010000011101001100;
		b = 32'b00000101011000110001000101111010;
		correct = 32'b10111000111010111111110100011011;
		#400 //-1.0539604e+31 * 1.0676699e-35 = -0.00011252818
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110010000001101010010101001111;
		b = 32'b00111010101111100101011100001101;
		correct = 32'b11101101010010000011100011110011;
		#400 //-2.6669336e+30 * 0.0014521793 = -3.8728656e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001011110001111110101111001110;
		b = 32'b11111110111010100011101011000001;
		correct = 32'b01001011001101101110101101101100;
		#400 //-7.700681e-32 * -1.5567221e+38 = 11987820.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110100100110111110100001111001;
		b = 32'b00011010100001001100101101010010;
		correct = 32'b10001111101000011011111101100011;
		#400 //-2.9040146e-07 * 5.49224e-23 = -1.5949545e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101111111101100111011111000011;
		b = 32'b10001100011001101011010000011100;
		correct = 32'b00111100110111100001110100000000;
		#400 //-1.5255619e+29 * -1.7772755e-31 = 0.027113438
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110001100000111101110011110010;
		b = 32'b11110110010100111011110001100111;
		correct = 32'b11101000010110100010000001001110;
		#400 //3.8377204e-09 * -1.0736288e+33 = -4.1202872e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111010010100100100101011010010;
		b = 32'b10011111010001100100000011010110;
		correct = 32'b01011010001000101101101100100001;
		#400 //-2.7297497e+35 * -4.1981762e-20 = 1.145997e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110001010110110110101110010;
		b = 32'b01110010110001100110110101000010;
		correct = 32'b01110001100001001101111111010000;
		#400 //0.16740969 * 7.860495e+30 = 1.315923e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000001000001111110011110011001;
		b = 32'b11101000111101110111100100000000;
		correct = 32'b00101010100000110110000010110001;
		#400 //-2.4961747e-38 * -9.3492526e+24 = 2.3337368e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101110101110000111111100100011;
		b = 32'b01001010101100101101101000000100;
		correct = 32'b00111010000000001110010110000101;
		#400 //8.389935e-11 * 5860610.0 = 0.00049170136
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001110011101010001011010000100;
		b = 32'b10000000101000000111100101110011;
		correct = 32'b10001111100110011010001001011000;
		#400 //1027973400.0 * -1.4737247e-38 = -1.5149497e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011101110010100110000000100011;
		b = 32'b11001011001010111011101100001101;
		correct = 32'b00101001100001111100001000010110;
		#400 //-5.3568358e-21 * -11254541.0 = 6.028873e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111101011101011100110111000111;
		b = 32'b00010110101000010101000111100100;
		correct = 32'b00010100100110101110010100001011;
		#400 //0.060010698 * 2.6062633e-25 = 1.5640368e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010000011010111000100100000001;
		b = 32'b11110011100010000101001001011100;
		correct = 32'b11000100011110101101100100011110;
		#400 //4.6451122e-29 * -2.1601038e+31 = -1003.39246
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000110100001100000100110010100;
		b = 32'b01000001011001110101101001001011;
		correct = 32'b01001000011100100100001111010110;
		#400 //17156.79 * 14.459544 = 248079.34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101001110111000001110110001000;
		b = 32'b11100011001011101010000011100110;
		correct = 32'b11001101100101100010011001101011;
		#400 //9.7750855e-14 * -3.2213274e+21 = -314887520.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100000000110010110001101110010;
		b = 32'b00111001100111001111000011101000;
		correct = 32'b10011010001111000001000111100011;
		#400 //-1.2992508e-19 * 0.00029934128 = -3.8891938e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010000010011100100001011010101;
		b = 32'b01000110111000001011000011110110;
		correct = 32'b00010111101101010000100100001111;
		#400 //4.0677822e-29 * 28760.48 = 1.1699138e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110101000011101110000000000101;
		b = 32'b10111011001101100010111111100001;
		correct = 32'b00110000110010110101101111111001;
		#400 //-5.3225114e-07 * -0.0027799534 = 1.4796334e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111100011011011001110101111111;
		b = 32'b00111100110101111111011100001111;
		correct = 32'b01111001110010000111010010010111;
		#400 //4.935075e+36 * 0.026362924 = 1.3010301e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100010000111010010100011011011;
		b = 32'b01000110001110110111001001101101;
		correct = 32'b00101000111001100010011000101110;
		#400 //2.1299096e-18 * 11996.606 = 2.5551687e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100101101001101111111100011001;
		b = 32'b01001111010001100110110101110000;
		correct = 32'b01110101100000010111000010110001;
		#400 //9.857732e+22 * 3329060900.0 = 3.281699e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000001110011011100010010111001;
		b = 32'b01010010011000000010100010000010;
		correct = 32'b10010100101101000010110010110001;
		#400 //-7.558739e-38 * 240688070000.0 = -1.8192983e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000110100011100111110001001100;
		b = 32'b00001011010110000100100111001111;
		correct = 32'b10010010011100001100001111101010;
		#400 //-18238.148 * 4.1655614e-32 = -7.597213e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100011101101111010110101011000;
		b = 32'b00110100111011000110101110001111;
		correct = 32'b01011001001010011010000011111001;
		#400 //6.77649e+21 * 4.4036685e-07 = 2984141400000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100011001001110110010101000010;
		b = 32'b01000111101111111010000101011010;
		correct = 32'b11101011011110101001110000011100;
		#400 //-3.0879027e+21 * 98114.7 = -3.0296866e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000001001101110110101100101000;
		b = 32'b11100010010011010011000000110101;
		correct = 32'b00100100000100110000001101011001;
		#400 //-3.3688672e-38 * -9.4626405e+20 = 3.187838e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110010111001110001000010010111;
		b = 32'b11000001101000111011011000111101;
		correct = 32'b01110101000100111100010000001101;
		#400 //-9.15342e+30 * -20.463984 = 1.8731543e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000000001001001010110010101011;
		b = 32'b10111100010010011001110011100100;
		correct = 32'b10111101000000011011000001111110;
		#400 //2.5730388 * -0.012305472 = -0.031662457
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011111000111001110101110010110;
		b = 32'b11110101000001110110110100100001;
		correct = 32'b11010100101001100000011001000001;
		#400 //3.3229157e-20 * -1.7167321e+32 = -5704556000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110011010011110010100011000010;
		b = 32'b10001000111100101011110001010011;
		correct = 32'b10111100110001000110110011101100;
		#400 //1.6412844e+31 * -1.460912e-33 = -0.02397772
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111001111001001100111001001;
		b = 32'b01110011001001101111001010011101;
		correct = 32'b11101010111101011111110011101011;
		#400 //-1.1241479e-05 * 1.322696e+31 = -1.486906e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010000000101010000011100100110;
		b = 32'b01011011000000101010010110101001;
		correct = 32'b10101011100110000001110000100011;
		#400 //-2.9390576e-29 * 3.6773892e+16 = -1.0808059e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010110000101000001101111100110;
		b = 32'b10000111101111000011101001010100;
		correct = 32'b00011110010110011100110001111000;
		#400 //-40711886000000.0 * -2.8321378e-34 = 1.15301675e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101011111010101110010111011001;
		b = 32'b10010101000001000100001011000010;
		correct = 32'b10000001011100101011011110001010;
		#400 //1.6690496e-12 * -2.670985e-26 = -4.4580063e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010011111010011010001110010011;
		b = 32'b01001011010000100010100010111100;
		correct = 32'b01011111101100010011001100100011;
		#400 //2006943400000.0 * 12724412.0 = 2.5537176e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010010101011110100111111000000;
		b = 32'b00111011100100110001110101100001;
		correct = 32'b01001110110010010111110111010011;
		#400 //376478630000.0 * 0.004489586 = 1690233200.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111001100110110101001100000000;
		b = 32'b10010001000000001101010101100101;
		correct = 32'b01001011000111000101010111110011;
		#400 //-1.0081118e+35 * -1.0163177e-28 = 10245619.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011011101010001001101011110101;
		b = 32'b00011010000111101000011010000000;
		correct = 32'b10110110010100001101000001110001;
		#400 //-9.491635e+16 * 3.2782282e-23 = -3.1115744e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110000011011101001001111100;
		b = 32'b10101100011111101001001110110111;
		correct = 32'b00100011000011010000100010101100;
		#400 //-2.1133155e-06 * -3.617757e-12 = 7.645462e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111101101001001111110111000001;
		b = 32'b10100010010010000010000111100011;
		correct = 32'b10100000100000001111110000010110;
		#400 //0.08056212 * -2.7122994e-18 = -2.185086e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100110011100111010111000010001;
		b = 32'b10100010001010001110100111110100;
		correct = 32'b00001001001000001100100011101101;
		#400 //-8.4543465e-16 * -2.28921e-18 = 1.9353774e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001000101101101000000001101111;
		b = 32'b11010001100111111001111011100000;
		correct = 32'b10011010111000111001011000010000;
		#400 //1.0983921e-33 * -85695660000.0 = -9.412744e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101010000100101111110101010010;
		b = 32'b01011111111010111101011100011101;
		correct = 32'b01001010100001110110101000001110;
		#400 //1.3055293e-13 * 3.3988167e+19 = 4437255.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001111100110111000101001000001;
		b = 32'b11010100001100011001000100011100;
		correct = 32'b00100100010101111100010110000011;
		#400 //-1.5337434e-29 * -3050575000000.0 = 4.6787992e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010010101010111011101110011;
		b = 32'b11101001011001011000010110111100;
		correct = 32'b01100100001111110110001101011110;
		#400 //-0.00081431045 * -1.7342222e+25 = 1.4121953e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010111000010001010001001101101;
		b = 32'b10101000010001101111010101111111;
		correct = 32'b10111111110101000110000101001111;
		#400 //150231200000000.0 * -1.1044441e-14 = -1.6592196
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001100010111010100010001110101;
		b = 32'b01011111011111110101000101000111;
		correct = 32'b10101100010111001010110101110001;
		#400 //-1.7045821e-31 * 1.8397564e+19 = -3.136016e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001101000000001011010101100010;
		b = 32'b01101111101000101100101111111011;
		correct = 32'b00111101001000111011001010101100;
		#400 //3.9661377e-31 * 1.0076634e+29 = 0.039965317
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110100101001100100110011100111;
		b = 32'b01010100110101101101001011111010;
		correct = 32'b11001010000010111000110101010111;
		#400 //-3.0975863e-07 * 7381301000000.0 = -2286421.8
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011101000011110001101111000011;
		b = 32'b01100000000100101110001100001000;
		correct = 32'b11111101101001000011100101111111;
		#400 //-6.4450314e+17 * 4.233725e+19 = -2.728649e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010000100110101100101011000011;
		b = 32'b00110110110100111000011111101011;
		correct = 32'b10000111111111111100111010011011;
		#400 //-6.1054694e-29 * 6.304113e-06 = -3.8489567e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011110010100111011100100001011;
		b = 32'b00111100101100111110100011101010;
		correct = 32'b01011011100101001100101100000100;
		#400 //3.8140593e+18 * 0.021961648 = 8.376303e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101101101101101010110000000001;
		b = 32'b01100001110000101101010110101110;
		correct = 32'b01010000000010110000011011010010;
		#400 //2.076739e-11 * 4.492582e+20 = 9329920000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001001111000100011100010010001;
		b = 32'b01000000101111110110100100001100;
		correct = 32'b10001011001010010010010100001000;
		#400 //-5.4460716e-33 * 5.981573 = -3.2576075e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110010011011111001000110011100;
		b = 32'b00101010011100011111100110011011;
		correct = 32'b11011101011000100111000110101010;
		#400 //-4.7451487e+30 * 2.1491699e-13 = -1.0198131e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010110110100000101111010100101;
		b = 32'b01011111001000100011001110001100;
		correct = 32'b01110110100001000000010111011001;
		#400 //114552460000000.0 * 1.1687839e+19 = 1.3388707e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110100100011110000101110101110;
		b = 32'b00110101011011110010001111101001;
		correct = 32'b10101010100001011001111111111000;
		#400 //-2.6644324e-07 * 8.9086694e-07 = -2.3736547e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011110111001011110000111110101;
		b = 32'b10110100000000100100010110011000;
		correct = 32'b11010011011010011111011001111010;
		#400 //8.282395e+18 * -1.2132512e-07 = -1004862600000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111000101100111100110100010010;
		b = 32'b10110001011110000001000101010100;
		correct = 32'b01101010101011100011101011010101;
		#400 //-2.917439e+34 * -3.60986e-09 = 1.0531546e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001100111011010011100000011010;
		b = 32'b00101000010100000000000101001100;
		correct = 32'b10110101110000001011111011001001;
		#400 //-124371150.0 * 1.1546601e-14 = -1.436064e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011000110000010111101000100110;
		b = 32'b11000101000101111011010010111111;
		correct = 32'b11011110011001010100111101001101;
		#400 //1701843000000000.0 * -2427.2966 = -4.1308776e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110101101001101010001001001;
		b = 32'b11100011100010001110111110000010;
		correct = 32'b01011010110000010111001111101010;
		#400 //-5.3891313e-06 * -5.052031e+21 = 2.722606e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011001110011001110010110011110;
		b = 32'b11010110001011100100000101110101;
		correct = 32'b01110000100010110111100001110101;
		#400 //-7209170000000000.0 * -47899040000000.0 = 3.4531232e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110010110000100110010000100000;
		b = 32'b00111000111101100001010000000100;
		correct = 32'b01101100001110101101101101101010;
		#400 //7.7006254e+30 * 0.00011733922 = 9.035854e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110010010011100100100110111;
		b = 32'b01010110010001111010001010110000;
		correct = 32'b11001101000111010101101110100110;
		#400 //-3.0068456e-06 * 54875388000000.0 = -165001820.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010000110011110000110010001010;
		b = 32'b10110111101001110011101011011000;
		correct = 32'b11001001000001110100000011000110;
		#400 //27789644000.0 * -1.9935353e-05 = -553996.4
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000000011110111011100011101001;
		b = 32'b01001010000000110110001001111001;
		correct = 32'b11001011000000010011000001110011;
		#400 //-3.933161 * 2152606.2 = -8466547.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000110110100111000101100100100;
		b = 32'b01000011100010011100100111001101;
		correct = 32'b10001010111000111011100001110000;
		#400 //-7.957383e-35 * 275.57657 = -2.1928683e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111101000000010011001001101111;
		b = 32'b11011001011101000000100111100000;
		correct = 32'b01010110111101100101001000011011;
		#400 //-0.031542238 * -4293172000000000.0 = 135416250000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101000100011111110101010111010;
		b = 32'b00110100011110001011100100100100;
		correct = 32'b00011101100010111101001101111001;
		#400 //1.5977986e-14 * 2.3164154e-07 = 3.701165e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110010110110001110101001001100;
		b = 32'b10101010101111100001111010001011;
		correct = 32'b01011110001000010001011111000110;
		#400 //-8.592897e+30 * -3.3771973e-13 = 2.901991e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011010101111001011111100101100;
		b = 32'b11110001101110101011011110011000;
		correct = 32'b01001101000010011010101001000011;
		#400 //-7.806383e-23 * -1.8491572e+30 = 144352300.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100111111111000100001010011111;
		b = 32'b01101110001100100001011100000101;
		correct = 32'b11010110101011110111110100000001;
		#400 //-7.001628e-15 * 1.377904e+28 = -96475710000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011011000000010010011011001111;
		b = 32'b11001100101100000011001011101001;
		correct = 32'b01101000001100011100100010111011;
		#400 //-3.6352942e+16 * -92378950.0 = 3.3582468e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101100000001010010000001011001;
		b = 32'b11001101000010011000011000100001;
		correct = 32'b01111001100011110000100000011111;
		#400 //-6.437596e+26 * -144204300.0 = 9.28329e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011001011111001111010101001000;
		b = 32'b10010001100010101100111111000111;
		correct = 32'b10101011100010010010100110001000;
		#400 //4450086500000000.0 * -2.1900614e-28 = -9.745963e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101110101000111011011110000010;
		b = 32'b11001111001100111110010011011000;
		correct = 32'b00111110011001100001011101010011;
		#400 //-7.4449794e-11 * -3018119200.0 = 0.22469835
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011010111001110000000001110110;
		b = 32'b11100111100000000000110100011100;
		correct = 32'b01000010111001110001100000011111;
		#400 //-9.5540105e-23 * -1.2094095e+24 = 115.54711
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011001011101010110100000110000;
		b = 32'b01000001101100101100101111000010;
		correct = 32'b11011011101010110110010111000101;
		#400 //-4317245300000000.0 * 22.349491 = -9.6488236e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000100000100010110001000001011;
		b = 32'b10110010001011100100001111000011;
		correct = 32'b00110110110001011110111000111110;
		#400 //-581.5319 * -1.014354e-08 = 5.8987926e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110001001110000010011111010000;
		b = 32'b10000111110110000011101011100101;
		correct = 32'b10111001100110111000101111110101;
		#400 //9.1189395e+29 * -3.2534683e-34 = -0.0002966818
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001001100101000000001100001000;
		b = 32'b11011001100110111000011011010111;
		correct = 32'b00100011101100111101011110010111;
		#400 //-3.5632555e-33 * -5472110000000000.0 = 1.9498525e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001100100011101010011010100001;
		b = 32'b11101101010110011111000100101100;
		correct = 32'b01111010011100101110001101000100;
		#400 //-74790150.0 * -4.215613e+27 = 3.1528633e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010011000100110010000111100010;
		b = 32'b00111010001110110100001001001000;
		correct = 32'b01001101110101110011111110110000;
		#400 //631928650000.0 * 0.00071433606 = 451409400.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110100111111111101011010100000;
		b = 32'b11101000101110110110000101000011;
		correct = 32'b11011110001110110100001011111010;
		#400 //4.7653612e-07 * -7.0790136e+24 = -3.3734056e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110011111010000011000101010100;
		b = 32'b00001011001111000000111101101101;
		correct = 32'b10111111101010101001001000110111;
		#400 //-3.67924e+31 * 3.6219088e-32 = -1.3325871
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011001110111110011010001101000;
		b = 32'b01111100001100011001000100010100;
		correct = 32'b01010110100110101101000110111010;
		#400 //2.3078826e-23 * 3.6879163e+36 = 85112780000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101001011100110111010111111101;
		b = 32'b11010000101010111001110101101101;
		correct = 32'b10111010101000110011010110000111;
		#400 //5.4059178e-14 * -23033768000.0 = -0.0012451865
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101100001101000001010010100110;
		b = 32'b11001010000010111101011111010100;
		correct = 32'b11110110110001001011111000010001;
		#400 //8.708166e+26 * -2291189.0 = -1.9952054e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001001010010011111111010001101;
		b = 32'b00100011101010111011111101111011;
		correct = 32'b10101101100001111000010000011110;
		#400 //-827368.8 * 1.8620952e-17 = -1.5406395e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000001010101101011111110001010;
		b = 32'b01010101100000101100100110100010;
		correct = 32'b01010111010110110110110011010001;
		#400 //13.421762 * 17975315000000.0 = 241260410000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011010100110101101001010010011;
		b = 32'b11010111011000010000010100011010;
		correct = 32'b01110010100010000001011000101001;
		#400 //-2.1789338e+16 * -247412030000000.0 = 5.390944e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101111100101000110010001100111;
		b = 32'b10101110010110001111100100000100;
		correct = 32'b11011110011110111000101000011110;
		#400 //9.185032e+28 * -4.9333884e-11 = -4.5313332e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110100000001000000100011100;
		b = 32'b11001111011000011111011001110000;
		correct = 32'b11001110011000101101101001011100;
		#400 //0.25098503 * -3791024000.0 = -951490300.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111111111100110010010001110011;
		b = 32'b00011101010100010010100101101100;
		correct = 32'b10011101110001101010100000011001;
		#400 //-1.8995498 * 2.7682334e-21 = -5.2583973e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100111001010111000111011010011;
		b = 32'b01010011101000010001010101111111;
		correct = 32'b01111011010101111110011001110101;
		#400 //8.101593e+23 * 1383700800000.0 = 1.12101805e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001010101001110000000000101100;
		b = 32'b11101001100111111101101110011001;
		correct = 32'b01110100110100001001000010111001;
		#400 //-5472278.0 * -2.4157028e+25 = 1.3219398e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011101111110100001011001100101;
		b = 32'b01001100111000010100001011000101;
		correct = 32'b00101011010111000000111011101001;
		#400 //6.6197604e-21 * 118101544.0 = 7.8180393e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101100010100010111001111000001;
		b = 32'b11101100101001100100001001110000;
		correct = 32'b11011001100010000000011101101011;
		#400 //2.9764943e-12 * -1.6079634e+27 = -4786094000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011010100000011111010101110101;
		b = 32'b01001001101110000001100111101011;
		correct = 32'b00100100101110101110101100101001;
		#400 //5.3749707e-23 * 1508157.4 = 8.106302e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000111000011000101011000110100;
		b = 32'b01001001000101110001100101001010;
		correct = 32'b10010000101001011010100101101011;
		#400 //-1.0557762e-34 * 618900.6 = -6.5342054e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110110010011010110110100100110;
		b = 32'b10001101100011111100100000010111;
		correct = 32'b11000100011001101100000100010000;
		#400 //1.0416354e+33 * -8.861225e-31 = -923.0166
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100111101110100100100111100000;
		b = 32'b01101101001010110010101000101110;
		correct = 32'b01010101011110010001110000010100;
		#400 //5.1705466e-15 * 3.310808e+27 = 17118687000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111101011101101101110100100100;
		b = 32'b00000111111100100000111011001011;
		correct = 32'b01000101111010010110101101010000;
		#400 //2.0508645e+37 * 3.6420808e-34 = 7469.414
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010111011011000110111101011001;
		b = 32'b01100010011011111001001110000001;
		correct = 32'b10111010010111010100010000101111;
		#400 //-7.6396253e-25 * 1.10485015e+21 = -0.0008440641
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000101101010011111000010110000;
		b = 32'b01001110111100101011101001000111;
		correct = 32'b10010101001000010010000100101110;
		#400 //-1.5981098e-35 * 2036147100.0 = -3.2539865e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010001111001111101110011011011;
		b = 32'b01111011001101001001110001011001;
		correct = 32'b11001101101000111001010011100101;
		#400 //-3.6581487e-28 * 9.3778454e+35 = -343055520.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100011101011001100111000011100;
		b = 32'b10100000101110001101001100010110;
		correct = 32'b00000100111110011000010101000010;
		#400 //-1.8735568e-17 * -3.1310497e-19 = 5.8661997e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010010101100110111000010010111;
		b = 32'b00010100000001111010000101011011;
		correct = 32'b10100111001111100010001011110010;
		#400 //-385344050000.0 * 6.84758e-27 = -2.638674e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101001011001001100011011100110;
		b = 32'b01000011011000011111011010100100;
		correct = 32'b00101101010010011110111100111010;
		#400 //5.0798687e-14 * 225.96344 = 1.1478646e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001100011000000000000001001101;
		b = 32'b10000011000101011011110110000110;
		correct = 32'b10010000000000110000011000000010;
		#400 //58720564.0 * -4.4004727e-37 = -2.5839823e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101010001010000110011010111011;
		b = 32'b11000001110110000101111110001001;
		correct = 32'b11101100100011100101010110000110;
		#400 //5.0896167e+25 * -27.046648 = -1.3765707e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111110011001111001110011111000;
		b = 32'b01111001111011010011010111100100;
		correct = 32'b11111000110101101001110100010011;
		#400 //-0.22618473 * 1.5395842e+35 = -3.4823043e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000011100000001010111101010001;
		b = 32'b11101011011111111100000100010011;
		correct = 32'b11101111100000001000111110101111;
		#400 //257.36966 * -3.0918785e+26 = -7.957557e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010000000001101010001001100001;
		b = 32'b11101000111001010100000001000111;
		correct = 32'b10111001011100010010001000011101;
		#400 //2.6551932e-29 * -8.660861e+24 = -0.00022996259
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100010000001010010011101101111;
		b = 32'b11001110111101011110001011010011;
		correct = 32'b11110001011111111100100101110000;
		#400 //6.140646e+20 * -2062641500.0 = -1.2665952e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101001001110100111110100010100;
		b = 32'b00001010111000100010001100110101;
		correct = 32'b10110100101001001011110000010001;
		#400 //-1.4090679e+25 * 2.1776252e-32 = -3.0684217e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101011000011110100111000011011;
		b = 32'b10101111101010000111000011100010;
		correct = 32'b01011011001111001001010011100101;
		#400 //-1.7324523e+26 * -3.063923e-10 = 5.3081007e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010111110010111110001110100000;
		b = 32'b10100101000111001011001100101101;
		correct = 32'b00111101011110011001101011010011;
		#400 //-448357000000000.0 * -1.359155e-16 = 0.060938668
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110111110010010101000010111;
		b = 32'b01010010000000101111010100010010;
		correct = 32'b01010001011111101110101111001101;
		#400 //0.48664925 * 140614340000.0 = 68429860000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001001100000001100010101100000;
		b = 32'b01011101000100000011100010101100;
		correct = 32'b01100111000100010001011100001111;
		#400 //1054892.0 * 6.495153e+17 = 6.851685e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100011000110101111101110110000;
		b = 32'b11010100101011011011100101001000;
		correct = 32'b01111000010100100101100010000011;
		#400 //-2.8589346e+21 * -5969103000000.0 = 1.7065275e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101111000111110101001001101001;
		b = 32'b10100101111111111010111010111100;
		correct = 32'b01010101100111110001111111010110;
		#400 //-4.9307744e+28 * -4.4353853e-16 = 21869885000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011011111100011011100011001011;
		b = 32'b10111110111101001011010001001101;
		correct = 32'b01011011011001110000111001100000;
		#400 //-1.360773e+17 * -0.4779381 = 6.5036525e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001111010011010111010100111111;
		b = 32'b01010100101010101100111001100001;
		correct = 32'b00100100100010010001010101111110;
		#400 //1.0129861e-29 * 5868855000000.0 = 5.945069e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011111011010000111110100010010;
		b = 32'b10111111000000010111010011011010;
		correct = 32'b00011110111010110010001001001001;
		#400 //-4.9231367e-20 * -0.50568926 = 2.4895773e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101110000010001010110100000100;
		b = 32'b10111110011110101011111001100101;
		correct = 32'b10101101000001011101111010011100;
		#400 //3.107649e-11 * -0.24486692 = -7.609604e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001000110010000000100100111100;
		b = 32'b11001001100101111100001111110110;
		correct = 32'b01010010111011010010110100100011;
		#400 //-409673.88 * -1243262.8 = 509332260000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111101000100011111000100001000;
		b = 32'b01110011101101110000111110111001;
		correct = 32'b11110001010100001011100010000111;
		#400 //-0.035630256 * 2.900724e+31 = -1.0335354e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100101000011011010110000101111;
		b = 32'b01000010000110010101101110100111;
		correct = 32'b11100111101010011011110101000001;
		#400 //-4.181437e+22 * 38.339504 = -1.6031421e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110111100000010000000100110001;
		b = 32'b01000000101100110001100101011000;
		correct = 32'b01111000101101001000000100110101;
		#400 //5.2330505e+33 * 5.5968437 = 2.9288565e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001001100111101101111100001011;
		b = 32'b10001001101001110001101100100110;
		correct = 32'b10010011110011110110100010110011;
		#400 //1301473.4 * -4.0229318e-33 = -5.2357388e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010111011111110001001111110011;
		b = 32'b00101101011000010000010011010011;
		correct = 32'b10000101011000000011010101010111;
		#400 //-8.2420123e-25 * 1.27908404e-11 = -1.05422264e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110101111100110111011011000000;
		b = 32'b11010110011100010111000000000110;
		correct = 32'b11001100111001011001110101010100;
		#400 //1.8139472e-06 * -66365860000000.0 = -120384160.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110110110101110011000000110000;
		b = 32'b11000100110110010101101101101011;
		correct = 32'b10111100001101101011010010110001;
		#400 //6.413109e-06 * -1738.8568 = -0.011151479
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100011101111000100011010011111;
		b = 32'b00110111000010100011001010000110;
		correct = 32'b10011011010010110100011001110100;
		#400 //-2.041291e-17 * 8.237204e-06 = -1.6814531e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010000010111100101101000100010;
		b = 32'b00110001000000101011000011100000;
		correct = 32'b11000001111000110000011011001100;
		#400 //-14921796000.0 * 1.9018032e-09 = -28.378319
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000100010110001010011110100100;
		b = 32'b11110001100111000001010101010000;
		correct = 32'b01110110100001000001100000110001;
		#400 //-866.6194 * -1.5457737e+30 = 1.3395974e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000001100101001100111001101;
		b = 32'b00100001011010011111100000100111;
		correct = 32'b10010010001000110011101100011100;
		#400 //-6.4974587e-10 * 7.92719e-19 = -5.150659e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001011100110010001011000101111;
		b = 32'b00110110011100101110000010001100;
		correct = 32'b01000010100100010011110101000000;
		#400 //20065374.0 * 3.6191514e-06 = 72.61963
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111100101011110011111000011000;
		b = 32'b01001010011001111101001100011111;
		correct = 32'b01000111100111101011000110001101;
		#400 //0.021391913 * 3798215.8 = 81251.1
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010001101010000101000000010110;
		b = 32'b11000111010110011111111000010111;
		correct = 32'b10011001100011110101001011110001;
		#400 //2.6555083e-28 * -55806.09 = -1.4819353e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010001101100101001000110100110;
		b = 32'b01101000101101111011000101111100;
		correct = 32'b00111011000000000010000111101011;
		#400 //2.817321e-28 * 6.9397366e+24 = 0.0019551467
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100111101101011011001101111010;
		b = 32'b01100110000000100010111001111110;
		correct = 32'b11001110001110001100110001000111;
		#400 //-5.043218e-15 * 1.5369132e+23 = -775098800.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101111111001010001100101100100;
		b = 32'b00100010001011011100001100000000;
		correct = 32'b10010010100110111000000010101011;
		#400 //-4.1672898e-10 * 2.3549104e-18 = -9.813594e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110100000000001110010110110000;
		b = 32'b01001010111100100001111010111100;
		correct = 32'b00111111011100111101000100110100;
		#400 //1.2004489e-07 * 7933790.0 = 0.95241094
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111011110101101011100001001010;
		b = 32'b01110001011010101111001010010111;
		correct = 32'b11101101110001010000111111101101;
		#400 //-0.0065527307 * 1.16340425e+30 = -7.623475e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110101101011110111100100011011;
		b = 32'b10011011010010100001111111011001;
		correct = 32'b01010001100010101000101101100100;
		#400 //-4.4487708e+32 * -1.6719339e-22 = 74380510000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000010001011011110011001111110;
		b = 32'b10000000100110001000010101110101;
		correct = 32'b00000011010011110011011100000110;
		#400 //-43.47509 * -1.4006871e-38 = 6.0894996e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110111000010001001101010111100;
		b = 32'b01100101110110101100000101110110;
		correct = 32'b01011101011010010111010111111111;
		#400 //8.142259e-06 * 1.2913058e+23 = 1.0514145e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110001111100110101100000001;
		b = 32'b10001110111001011110100101111100;
		correct = 32'b00000101101010110000001101100100;
		#400 //-2.837449e-06 * -5.6677696e-30 = 1.6082008e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011110001100000011101111011111;
		b = 32'b10001011010100110010110100010010;
		correct = 32'b10101010000100010110000001100000;
		#400 //3.1747472e+18 * -4.067103e-32 = -1.2912024e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010111001001111101000101100000;
		b = 32'b11110101111111010110010011001101;
		correct = 32'b01001101101001100001110000000000;
		#400 //-5.422488e-25 * -6.424295e+32 = 348356600.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110000110101010011000011011001;
		b = 32'b00110010011010001110101010111101;
		correct = 32'b00100011110000011111011111000001;
		#400 //1.5511673e-09 * 1.3557551e-08 = 2.103003e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101101000111001010110101100110;
		b = 32'b11011011000000111101001100100111;
		correct = 32'b11001000101000010101101111101100;
		#400 //8.9060755e-12 * -3.7105386e+16 = -330463.38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011010110100111101111110110100;
		b = 32'b01101100110101110100010010000110;
		correct = 32'b11001000001100100010100110010110;
		#400 //-8.7628967e-23 * 2.0819412e+27 = -182438.34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100000010111001110100101000100;
		b = 32'b10100000100111100011001100100111;
		correct = 32'b10000001100010001000010000011100;
		#400 //1.8711906e-19 * -2.680009e-19 = -5.014808e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011110100011010110011110111111;
		b = 32'b11000100110110100011000010110100;
		correct = 32'b11100011111100010000101001111111;
		#400 //5.0946613e+18 * -1745.522 = -8.8928433e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101010111011110101010010010100;
		b = 32'b00110110000110101110111010011100;
		correct = 32'b11100001100100001101011111110100;
		#400 //-1.4466634e+26 * 2.3086677e-06 = -3.3398653e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100010011011110000111001001011;
		b = 32'b10111100011110011110010101001101;
		correct = 32'b10011111011010010101101100000111;
		#400 //3.2398107e-18 * -0.0152524235 = -4.9414965e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111101011010111011011001101101;
		b = 32'b11001001101001100010100011010110;
		correct = 32'b11000111100110001111110111100100;
		#400 //0.05754702 * -1361178.8 = -78331.78
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001101000101100011110101001011;
		b = 32'b01011001010111011001110100001010;
		correct = 32'b01100111000000100000111100010011;
		#400 //157537460.0 * 3898664800000000.0 = 6.141857e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011010101100110000000000110011;
		b = 32'b11010111110001001111001101101101;
		correct = 32'b10110011000010011011011001011100;
		#400 //7.4032987e-23 * -433099570000000.0 = -3.2063653e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000011010101011010100111111111;
		b = 32'b11100001110011101111011111001011;
		correct = 32'b01100101101011001011110110011100;
		#400 //-213.66405 * -4.7723558e+20 = 1.0196809e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101000011111101100110010010011;
		b = 32'b01011001011011111001101000111011;
		correct = 32'b01000010011011100111101001111111;
		#400 //1.4144192e-14 * 4215131000000000.0 = 59.619625
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011110110000001111001101011;
		b = 32'b11101011001100010000111011110111;
		correct = 32'b01110111100101010111100110101010;
		#400 //-28327126.0 * -2.1405054e+26 = 6.0634365e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100111001100111110101001000;
		b = 32'b00011001100010110110011011110001;
		correct = 32'b00011110111110110000010101101010;
		#400 //1843.915 * 1.4413841e-23 = 2.6577898e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011101011111000100011111111100;
		b = 32'b00010000110110101100001110101000;
		correct = 32'b00101110110101111001011000011101;
		#400 //1.1361735e+18 * 8.6287295e-29 = 9.8037335e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100100111110011101011110001101;
		b = 32'b01110110110101011111111010001110;
		correct = 32'b11011100010100001101100011000111;
		#400 //-1.08351694e-16 * 2.1701606e+33 = -2.3514058e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011011111011110000101111011110;
		b = 32'b10101001011101100100000100111101;
		correct = 32'b00000101111001011111001001010010;
		#400 //-3.9546902e-22 * -5.4679558e-14 = 2.1624071e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001010101000001010000011011011;
		b = 32'b00010001110010011100100101111110;
		correct = 32'b10011100111111010011100101110011;
		#400 //-5263469.5 * 3.1836388e-28 = -1.6756986e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011011110101000000111010100110;
		b = 32'b10101010100111001100010000111001;
		correct = 32'b10000111000000011101101101111000;
		#400 //3.5081924e-22 * -2.7847324e-13 = -9.769377e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000110110110000010000011101110;
		b = 32'b11101100100000000000111000101001;
		correct = 32'b10110011110110000011100011010111;
		#400 //8.1298555e-35 * -1.238475e+27 = -1.0068623e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011101101111011010001010001;
		b = 32'b10110111101000111010110110110001;
		correct = 32'b01000011111010101110100011100111;
		#400 //-24078498.0 * -1.9511996e-05 = 469.81955
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000010010111001111111010000100;
		b = 32'b10010101111000001000101111001011;
		correct = 32'b10011000110000011101011101100001;
		#400 //55.24855 * -9.0693434e-26 = -5.0106808e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101101000101110100101001111011;
		b = 32'b01101100101011010010011101111000;
		correct = 32'b01011010010011001010100101010001;
		#400 //8.599894e-12 * 1.6746444e+27 = 1.4401765e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100111010011111110110001010111;
		b = 32'b00101111001110101100110010001100;
		correct = 32'b00010111000101111011011111011001;
		#400 //2.885514e-15 * 1.6989271e-10 = 4.902278e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100000010011011111100001010001;
		b = 32'b11110110110001010111001101000001;
		correct = 32'b11010111100111101101110011010001;
		#400 //1.7446336e-19 * -2.002383e+33 = -349342470000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111001010011110001000001101100;
		b = 32'b11001101011010010000111111010010;
		correct = 32'b11000111001111001000001010111110;
		#400 //0.00019747176 * -244383000.0 = -48258.742
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100100101001001110111111110110;
		b = 32'b00001010000100100100001010001110;
		correct = 32'b10101111001111000111011101110111;
		#400 //-2.4340456e+22 * 7.042162e-33 = -1.7140943e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001011110101101010000010101011;
		b = 32'b11000001010011101011101111001101;
		correct = 32'b11001101101011010101001010111101;
		#400 //28131670.0 * -12.92085 = -363485100.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001000111000011001011001100101;
		b = 32'b10101111001111111000001100111101;
		correct = 32'b00111000101010001100001011011011;
		#400 //-462003.16 * -1.7417974e-10 = 8.047159e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101011010011010101010001101011;
		b = 32'b00010111100101011011110001000100;
		correct = 32'b11000011011100000011001001000110;
		#400 //-2.4822845e+26 * 9.676424e-25 = -240.19638
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001001111111110111101000111001;
		b = 32'b11100000001110101101001000000010;
		correct = 32'b00101010101110100111000001100010;
		#400 //-6.1503955e-33 * -5.3847298e+19 = 3.3118218e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000111010010110010011011001;
		b = 32'b10011011001111111110011111111001;
		correct = 32'b00001100101011101111010110111011;
		#400 //-1.6981644e-09 * -1.5874104e-22 = 2.6956838e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000110001001101011111001000000;
		b = 32'b01000011001111111000010010101100;
		correct = 32'b00001001111110010111110010111000;
		#400 //3.1360904e-35 * 191.51825 = 6.0061854e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101101000011101011100100010111;
		b = 32'b00000100100101001111001010101110;
		correct = 32'b00110010001001100001010010011011;
		#400 //2.7606645e+27 * 3.50175e-36 = 9.667157e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000011001010111111000010110010;
		b = 32'b00100110011111111111010000101111;
		correct = 32'b10101010001010111110100011000010;
		#400 //-171.94022 * 8.880183e-16 = -1.5268605e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011000100100001110110101011100;
		b = 32'b00011010110011101001011011100101;
		correct = 32'b10110011111010011110100011011010;
		#400 //-1274793000000000.0 * 8.5443386e-23 = -1.08922634e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001111011001101010101111010101;
		b = 32'b11001100001011111011000100001110;
		correct = 32'b01011100000111100100111100000000;
		#400 //-3870020900.0 * -46056504.0 = 1.7823963e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000101101001000101101111110000;
		b = 32'b01010010010010111001100110100000;
		correct = 32'b11011000100000101011011110001001;
		#400 //-5259.492 * 218613940000.0 = -1149798300000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011101010000001100001010010110;
		b = 32'b11000110001001100110010001010101;
		correct = 32'b00100011111110101001001101110011;
		#400 //-2.5511587e-21 * -10649.083 = 2.7167501e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111001111101001101110100011110;
		b = 32'b01011000010001010001001110111011;
		correct = 32'b01010010101111001000000100000111;
		#400 //0.00046704052 * 866754100000000.0 = 404809300000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001010110101000010011011011011;
		b = 32'b01100011101101111110101100000001;
		correct = 32'b00101111000110000110101010000111;
		#400 //2.0429473e-32 * 6.785376e+21 = 1.3862166e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001110011000111011111111101101;
		b = 32'b01101011111000110111101111010101;
		correct = 32'b11111010110010100110000101011010;
		#400 //-955251500.0 * 5.500219e+26 = -5.2540924e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111001000110010010001010001011;
		b = 32'b01110111010100110100110010000010;
		correct = 32'b01110000111111001100101001111001;
		#400 //0.00014604085 * 4.28565e+33 = 6.2587998e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010010111011100110111001010000;
		b = 32'b00110000111001101100101111110111;
		correct = 32'b00000100010101101111010100010011;
		#400 //1.5047106e-27 * 1.6792673e-09 = 2.5268112e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001011011010110000111001111100;
		b = 32'b11110000101001000101111001010010;
		correct = 32'b10111100100101101110101111100010;
		#400 //4.527025e-32 * -4.0695654e+29 = -0.018423025
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001111100101001001010001010100;
		b = 32'b01001101001100010000001101100101;
		correct = 32'b01011101010011010111100100001101;
		#400 //4985497600.0 * 185611860.0 = 9.253675e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000010010001001101101010101000;
		b = 32'b11100000000100010111001000111011;
		correct = 32'b11100010110111111010111101100000;
		#400 //49.21353 * -4.1922017e+19 = -2.0631305e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010000111100100100110101110011;
		b = 32'b10001111000011000111100100010010;
		correct = 32'b00100000100001001111010011110011;
		#400 //-32521296000.0 * -6.92585e-30 = 2.2523764e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100101000011100000100110101000;
		b = 32'b10101110011011001000001001000100;
		correct = 32'b01010100000000110011100100101110;
		#400 //-4.1922135e+22 * -5.3775887e-11 = 2254400000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010010110111101111111110011110;
		b = 32'b10111100100100111001100000111011;
		correct = 32'b01010000000000001001000101100011;
		#400 //-478885640000.0 * -0.018016925 = 8628047000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011001001011100100010111100111;
		b = 32'b00000011001100110100110110111110;
		correct = 32'b10011100111101000001111110011010;
		#400 //-3065844000000000.0 * 5.2692616e-37 = -1.6154734e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011010101111000100100011011111;
		b = 32'b01001110010110001001110001000111;
		correct = 32'b01101001100111110101000001101101;
		#400 //2.649871e+16 * 908530100.0 = 2.4074876e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001001001101101010001000000011;
		b = 32'b10100010110011110111110110000101;
		correct = 32'b10101100100101000000011010001100;
		#400 //748064.2 * -5.624036e-18 = -4.20714e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011101001010111001101001001111;
		b = 32'b11101100100000100101111110011101;
		correct = 32'b11001010001011101100100011100111;
		#400 //2.2711437e-21 * -1.260895e+27 = -2863673.8
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111100001110010001011101110100;
		b = 32'b10000001101010101011101001101111;
		correct = 32'b00111110011101101110000010111101;
		#400 //-3.8442024e+36 * -6.2715656e-38 = 0.24109168
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101100000110110001111010011101;
		b = 32'b11001101101000010100101000100001;
		correct = 32'b11111010010000110111011001010111;
		#400 //7.501123e+26 * -338248740.0 = -2.5372453e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110000011100110111111100111100;
		b = 32'b01001000100000010100010001110001;
		correct = 32'b01111001011101011110100001101101;
		#400 //3.014347e+29 * 264739.53 = 7.980168e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001000101001100111011110100001;
		b = 32'b11000011011110110111000100100110;
		correct = 32'b10001100101000111000000011011110;
		#400 //1.0018886e-33 * -251.44199 = -2.5191686e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001001010110010110011111011001;
		b = 32'b01101101110010010001011100011100;
		correct = 32'b00110111101010101100011000101001;
		#400 //2.6169254e-33 * 7.779303e+27 = 2.0357855e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000110001001101001000111111000;
		b = 32'b01101001001000110110000101100100;
		correct = 32'b00101111110101001001110010011111;
		#400 //3.132837e-35 * 1.2344676e+25 = 3.867386e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000001001001111111001000000011;
		b = 32'b01000100001000111010101111000111;
		correct = 32'b10000101110101101011111110010010;
		#400 //-3.084669e-38 * 654.684 = -2.0194835e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011111100010101011001001000001;
		b = 32'b10000011000000111110010001100100;
		correct = 32'b10100011000011101110100111101000;
		#400 //1.9988244e+19 * -3.875962e-37 = -7.747367e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110001110000001011000001001111;
		b = 32'b00011100101101101000101100111101;
		correct = 32'b10001111000010010110011000100110;
		#400 //-5.6079794e-09 * 1.2079742e-21 = -6.7742946e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100011101100100010110010110000;
		b = 32'b01011111001010110110010000000001;
		correct = 32'b11000011011011101001001011100111;
		#400 //-1.9317725e-17 * 1.2349997e+19 = -238.57384
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110010001010001101000110111001;
		b = 32'b00100101101110100100101011101101;
		correct = 32'b01011000011101011011001110010011;
		#400 //3.3438093e+30 * 3.2316628e-16 = 1080606460000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010001101111100101011110110000;
		b = 32'b00110110111001011000111110010010;
		correct = 32'b11001001001010101010111100110000;
		#400 //-102189370000.0 * 6.8414456e-06 = -699123.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001011110110000101001001110101;
		b = 32'b10111010010000011111011110000010;
		correct = 32'b10000110101000111110011101010000;
		#400 //8.332424e-32 * -0.0007399247 = -6.165367e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011100100000001111010000000101;
		b = 32'b10101111011110110111100101001010;
		correct = 32'b01001100011111010101100010110011;
		#400 //-2.903768e+17 * -2.2871408e-10 = 66413260.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111101000000110101110111110010;
		b = 32'b01000011100011011101101010000010;
		correct = 32'b11000001000100011001010110111110;
		#400 //-0.032072015 * 283.7071 = -9.099058
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011100111101001001101101110110;
		b = 32'b01001101100110010101111011011001;
		correct = 32'b10101011000100101000101110001010;
		#400 //-1.6186751e-21 * 321641250.0 = -5.206327e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110011101011000101000000111000;
		b = 32'b00000000111111011110101110101101;
		correct = 32'b10110101001010101110100111101001;
		#400 //-2.730414e+31 * 2.3318925e-38 = -6.367032e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111110000110000000110101100100;
		b = 32'b10101100101001010011000110110001;
		correct = 32'b01101011010001000011110001001010;
		#400 //-5.0528046e+37 * -4.695099e-12 = 2.3723417e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001010010011001010011000101011;
		b = 32'b00010110101001001111111000111001;
		correct = 32'b00100001100000111110010110101110;
		#400 //3352970.8 * 2.6656066e-25 = 8.937701e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000001000110011101101110011100;
		b = 32'b01101100000111000001110011001011;
		correct = 32'b11101101101110111010011001000010;
		#400 //-9.616116 * 7.549136e+26 = -7.259336e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110110100010010101010110000;
		b = 32'b10110101101111011100000001000110;
		correct = 32'b10110101000110110000100110011101;
		#400 //0.4085288 * -1.4137556e-06 = -5.775599e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011100100001110001011111100011;
		b = 32'b10110001101100101110111001101010;
		correct = 32'b10001110101111001101100011011000;
		#400 //8.939725e-22 * -5.2075864e-09 = -4.655439e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010100000000101010000101100100;
		b = 32'b11001011001100101100110011011000;
		correct = 32'b11011111101101100111100101111101;
		#400 //2244213700000.0 * -11717848.0 = -2.6297356e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101011000010110100111001010101;
		b = 32'b01001110010000111010100000110101;
		correct = 32'b01111001110101001111000001100110;
		#400 //1.684106e+26 * 820645200.0 = 1.3820535e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000101001001000111011011111111;
		b = 32'b11000100111000000111101000100010;
		correct = 32'b10001010100100000011011010010110;
		#400 //7.733099e-36 * -1795.8167 = -1.3887229e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100111000000010110010000010110;
		b = 32'b11111111110000011011011100010011;
		correct = 32'b11111111110000011011011100010011;
		#400 //-1.7956603e-15 * nan = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001110000011001010100011110100;
		b = 32'b01000000000001100100000100111001;
		correct = 32'b01001110100100111000100010001100;
		#400 //589970700.0 * 2.0977309 = 1237599700.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011000101100001010110000010101;
		b = 32'b01111111110100001101111110101101;
		correct = 32'b01111111110100001101111110101101;
		#400 //-4.5668692e-24 * nan = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100110110101010000110110000000;
		b = 32'b11001011000010011101110101110110;
		correct = 32'b01110010011001010111100100010001;
		#400 //-5.0305655e+23 * -9035126.0 = 4.5451794e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001100011011110010011000110110;
		b = 32'b10011000101111111011111001000010;
		correct = 32'b10100101101100110001111100111110;
		#400 //62691544.0 * -4.9564454e-24 = -3.107272e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101011110000111011000111000110;
		b = 32'b00110101001111010111000011100100;
		correct = 32'b00100001100100001101000010001011;
		#400 //1.3904925e-12 * 7.0572264e-07 = 9.81302e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111111101010101011100010110010;
		b = 32'b11001100101110010011111111110111;
		correct = 32'b01001100111101110001010001000010;
		#400 //-1.3337615 * -97124280.0 = 129540620.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110101110100110110001001000111;
		b = 32'b00001100100001111001010011100100;
		correct = 32'b11000010110111111110011110001001;
		#400 //-5.3592184e+32 * 2.0889654e-31 = -111.95222
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000010010110010010011010010111;
		b = 32'b01011100000101111110101001010011;
		correct = 32'b01011111000000001101110010000111;
		#400 //54.287685 * 1.7104145e+17 = 9.285445e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100010001000110000111000000001;
		b = 32'b01101100111011011001000111111101;
		correct = 32'b11001111100101110101000011110011;
		#400 //-2.2098033e-18 * 2.2976386e+27 = -5077329400.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011111001000010010000111000000;
		b = 32'b10111010110100000010101011011101;
		correct = 32'b01011010100000110000011001100111;
		#400 //-1.1610772e+19 * -0.0015881915 = 1.844013e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101100000110011001110111101011;
		b = 32'b00111111111100111000100100011111;
		correct = 32'b00101100100100100010001100101110;
		#400 //2.183027e-12 * 1.9026221 = 4.1534753e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100101100100100110111101100010;
		b = 32'b10110110000000001110010011101101;
		correct = 32'b10011100000100110111010101001000;
		#400 //2.540244e-16 * -1.9206739e-06 = -4.87898e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110010110000011101011000111001;
		b = 32'b10111110100011000011100010001010;
		correct = 32'b01110001110101000101011111101101;
		#400 //-7.678667e+30 * -0.27386886 = 2.1029478e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010110101111111111000100110101;
		b = 32'b11010101101110011000111111010001;
		correct = 32'b01101101000010110010000100100100;
		#400 //-105521350000000.0 * -25503417000000.0 = 2.691155e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101100001011010101111000110001;
		b = 32'b11011100010011011110010010111111;
		correct = 32'b01001001000010110110111101010110;
		#400 //-2.4637065e-12 * -2.3181552e+17 = 571125.4
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001000001110000011001110011110;
		b = 32'b00100001110001001101110011010000;
		correct = 32'b10101010100011011010011001100111;
		#400 //-188622.47 * 1.3339925e-18 = -2.5162096e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100101010101101001111101010001;
		b = 32'b01010001000111010001010010011111;
		correct = 32'b00110111000000111011000011111110;
		#400 //1.861552e-16 * 42165990000.0 = 7.849418e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001010111000100110001101100111;
		b = 32'b01000111111001000010010111010000;
		correct = 32'b01010011010010011100000111111000;
		#400 //7418291.5 * 116811.625 = 866542700000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000111011011000011010011111110;
		b = 32'b10111100010111100010101001101011;
		correct = 32'b00000100010011001111110100011000;
		#400 //-1.777024e-34 * -0.013559918 = 2.40963e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101000101000001011000110001111;
		b = 32'b11100000111010111010011100101010;
		correct = 32'b01001010000100111110101111101100;
		#400 //-1.7840572e-14 * -1.358447e+20 = 2423547.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001110100101011010010100010010;
		b = 32'b01011101010010001100101001101101;
		correct = 32'b11101100011010101011111010010100;
		#400 //-1255311600.0 * 9.0428104e+17 = -1.1351545e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100110000100000011111010111110;
		b = 32'b11011111100100011111010111101111;
		correct = 32'b11000110001001000111110000111001;
		#400 //5.004507e-16 * -2.103515e+19 = -10527.056
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100011010011100101001011011101;
		b = 32'b11111100001110100110001010010001;
		correct = 32'b11100000000101100011011110100101;
		#400 //1.1184829e-17 * -3.8710655e+36 = -4.3297207e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111100000000110000110010001010;
		b = 32'b01001110000101111101100111110000;
		correct = 32'b01001010100110110111011111101100;
		#400 //0.007998595 * 636910600.0 = 5094390.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100011000111010100101111010001;
		b = 32'b00111100111000010001110000110000;
		correct = 32'b01100000100010100101000011110100;
		#400 //2.901602e+21 * 0.027479261 = 7.973387e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010100100000000100111110010;
		b = 32'b01000100011110100011110101111011;
		correct = 32'b10111111100011001100110001001110;
		#400 //-0.0010989292 * 1000.96063 = -1.0999849
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100111111001011110010101000010;
		b = 32'b00110010100011000101111111100100;
		correct = 32'b10011010111111000001111011111010;
		#400 //-6.380883e-15 * 1.6341751e-08 = -1.042748e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010100010011011100100110000011;
		b = 32'b00111100010111101010010001100001;
		correct = 32'b01010001001100101111100011100011;
		#400 //3535396400000.0 * 0.013588996 = 48042488000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000110000011011101100000110110;
		b = 32'b11001011100101101010100001101110;
		correct = 32'b01010010001001101111010000000101;
		#400 //-9078.053 * -19747036.0 = 179264630000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000010110010100000010011011011;
		b = 32'b01100010010100110110101101001011;
		correct = 32'b01100101101001101101011010101100;
		#400 //101.00948 * 9.749986e+20 = 9.84841e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001110101000101001110011111001;
		b = 32'b11011100111001000101101011001001;
		correct = 32'b10101100000100010000110101111001;
		#400 //4.0087242e-30 * -5.142089e+17 = -2.0613218e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101101001000001111101001011111;
		b = 32'b10100111100110110001111110100101;
		correct = 32'b11010101010000110001011011111011;
		#400 //3.1137676e+27 * -4.305545e-15 = -13406467000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000101010101101010010010011000;
		b = 32'b01100110111101100010011010100100;
		correct = 32'b11101100110011100110001010010000;
		#400 //-3434.287 * 5.8120747e+23 = -1.9960333e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011011000001101001111010101010;
		b = 32'b01000110101001001001001011001101;
		correct = 32'b10100010001011010001010110101110;
		#400 //-1.1135487e-22 * 21065.4 = -2.345735e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101001100000011110110010010110;
		b = 32'b10110000011100000010110010100101;
		correct = 32'b00011010011100111100100011101010;
		#400 //-5.769792e-14 * -8.7374935e-10 = 5.041352e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111111000000110001100011111110;
		b = 32'b01000001001001111011010000010010;
		correct = 32'b01000000101010111100001100001001;
		#400 //0.5121001 * 10.4814625 = 5.367558
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100110010101001111011100000100;
		b = 32'b11010010111010111001100101100100;
		correct = 32'b11111001110000111111111001011011;
		#400 //2.5142458e+23 * -505945400000.0 = -1.272071e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111110111001111000110111101101;
		b = 32'b01101111010111101001111100100001;
		correct = 32'b11101110110010010101110100000011;
		#400 //-0.45225468 * 6.8898047e+28 = -3.1159466e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011101001101100101110101000110;
		b = 32'b00000011000011100101010010010101;
		correct = 32'b10100000110010101100011111111011;
		#400 //-8.21296e+17 * 4.1827145e-37 = -3.4352467e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001010010100100001100001001010;
		b = 32'b11101000101001010101011100010001;
		correct = 32'b10110011100001111011000100011100;
		#400 //1.01157005e-32 * -6.2463725e+24 = -6.3186434e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101010111000110100001100100001;
		b = 32'b11001001110000010111010000000011;
		correct = 32'b01110101001010111011110010011001;
		#400 //-1.3737158e+26 * -1584768.4 = 2.1770214e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110101001010111000110100000000;
		b = 32'b10001001110011001000110001010000;
		correct = 32'b10111111100010010001001001100011;
		#400 //2.1746645e+32 * -4.9243163e-33 = -1.0708736
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111011000000011001110100010000;
		b = 32'b10110110111001011111110001011011;
		correct = 32'b00110010011010001110001010001000;
		#400 //-0.0019777454 * -6.85411e-06 = 1.3555685e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101101010000101011001111000100;
		b = 32'b11001110111111100101110000001000;
		correct = 32'b11111100110000010111010001011011;
		#400 //3.7660885e+27 * -2133722100.0 = -8.035786e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100001011001111001111011101001;
		b = 32'b01011100000100100001011011101000;
		correct = 32'b11111110000001000010110101011010;
		#400 //-2.6704054e+20 * 1.6448213e+17 = -4.3923394e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011000010000100100010010010000;
		b = 32'b10111001111011011110101011111101;
		correct = 32'b11010010101101001000101111001100;
		#400 //854398900000000.0 * -0.00045379243 = -387719760000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010011101000010010001010001101;
		b = 32'b11010111111000111100000011111111;
		correct = 32'b11101100000011110101101100011101;
		#400 //1384138800000.0 * -500836100000000.0 = -6.9322665e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010101110001011001110001001110;
		b = 32'b00111100001011011011111111100100;
		correct = 32'b10010010100001100001111011000000;
		#400 //-7.981427e-26 * 0.010604832 = -8.464169e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001100101011111111001111100101;
		b = 32'b01001110100011010000110111010000;
		correct = 32'b00011011110000011110010110100111;
		#400 //2.7109808e-31 * 1183246300.0 = 3.207758e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100011111101000110100111100111;
		b = 32'b00101000000110111011110011010001;
		correct = 32'b10001100100101001011000001100100;
		#400 //-2.6499384e-17 * 8.6451715e-15 = -2.2909172e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001011111010111011001110101110;
		b = 32'b10111010000101010111110011110111;
		correct = 32'b10000110100010011010001010100011;
		#400 //9.078906e-32 * -0.000570252 = -5.1772646e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011110110010001000000111010000;
		b = 32'b00000010100011111111101000101010;
		correct = 32'b00100001111000011000100011100110;
		#400 //7.224029e+18 * 2.1155549e-37 = 1.528283e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101101111110010100000001100011;
		b = 32'b11010000101001011101000111101000;
		correct = 32'b01111111001000010111001011011111;
		#400 //-9.642451e+27 * -22255976000.0 = 2.1460215e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001111011110100100100100101011;
		b = 32'b00110101111010111001101001010111;
		correct = 32'b01000101111001100101100000010000;
		#400 //4199099100.0 * 1.7553783e-06 = 7371.008
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010010111100010100000001111010;
		b = 32'b11011111101100000111111110100000;
		correct = 32'b10110011001001100101010010011010;
		#400 //1.5225133e-27 * -2.543612e+19 = -3.872683e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000101011000100011010001011110;
		b = 32'b01111111000010010110001000110110;
		correct = 32'b11000100111100101100100110011100;
		#400 //-1.0636087e-35 * 1.8261418e+38 = -1942.3003
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111101000001001111100101111100;
		b = 32'b01100000111101101011111011001101;
		correct = 32'b01011110100000000010101011011001;
		#400 //0.03246449 * 1.4223899e+20 = 4.6177163e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000001011110010100100000111111;
		b = 32'b01111011010101101110001100111111;
		correct = 32'b10111101010100010011111110101101;
		#400 //-4.578591e-38 * 1.1157606e+36 = -0.051086117
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011111000111100111101000001101;
		b = 32'b00111010000110001011110001010010;
		correct = 32'b10011001101111010001101000011000;
		#400 //-3.355876e-20 * 0.0005826402 = -1.9552681e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000111011011101110000110110111;
		b = 32'b01001101110001111010010001111101;
		correct = 32'b10010101101110100100101011110010;
		#400 //-1.7971462e-34 * 418680740.0 = -7.5243045e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110110111001000111101101000111;
		b = 32'b01100100011001111010000000111110;
		correct = 32'b01011011110011101011101001000001;
		#400 //6.809281e-06 * 1.7090978e+22 = 1.1637727e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001101110011011100111000111100;
		b = 32'b10000100010100011101111100101101;
		correct = 32'b10010010101010001011100011001010;
		#400 //431605630.0 * -2.467031e-36 = -1.0647845e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000000000111101111011101101011;
		b = 32'b01101101000111101111110011110100;
		correct = 32'b10101101000110011101101001101001;
		#400 //-2.843822e-39 * 3.075277e+27 = -8.74554e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111100000100010110100100100000;
		b = 32'b11010001000100011101011000110010;
		correct = 32'b01001101101001011010110001101011;
		#400 //-0.008875161 * -39147740000.0 = 347442530.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001111100111111101101001001111;
		b = 32'b01011010101010000101001011100111;
		correct = 32'b00101010110100100011011000010000;
		#400 //1.57627e-29 * 2.3689474e+16 = 3.7341007e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011000100001100110111101101001;
		b = 32'b00110000011010000111111000011010;
		correct = 32'b10001001011101000010111001011111;
		#400 //-3.4750684e-24 * 8.458031e-10 = -2.9392235e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110011110010100010001010000011;
		b = 32'b11111001100101101101101000000101;
		correct = 32'b01101101111011100011100010111100;
		#400 //-9.412636e-08 * -9.790831e+34 = 9.2157525e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101110100111001011110010000011;
		b = 32'b11001101011101010101001010011110;
		correct = 32'b11111100100101100011001011111110;
		#400 //2.425378e+28 * -257239520.0 = -6.23903e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011000101100101011111000001111;
		b = 32'b01100100011111010110111101001100;
		correct = 32'b01111101101100001111001110001010;
		#400 //1572234900000000.0 * 1.8700184e+22 = 2.9401082e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111110111011011011110101011111;
		b = 32'b10011100011111011000111100101101;
		correct = 32'b11011011111010110111100100011101;
		#400 //1.5800515e+38 * -8.389573e-22 = -1.3255957e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011001111000011001001010110111;
		b = 32'b10110001001000111110101111010111;
		correct = 32'b00001011100100000111000000111010;
		#400 //-2.3323712e-23 * -2.3853681e-09 = 5.563564e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110011010010011001010111001001;
		b = 32'b10110101110110110011011110111101;
		correct = 32'b11101001101011001001111100000111;
		#400 //1.5971217e+31 * -1.6332993e-06 = -2.6085778e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000111101010101111110010110100;
		b = 32'b10110010001101110110000110100000;
		correct = 32'b00111010011101001111011110110011;
		#400 //-87545.41 * -1.0674199e-08 = 0.00093447714
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100100100111010111001001010011;
		b = 32'b10011110000111101010011010110110;
		correct = 32'b10000011010000110010011000101111;
		#400 //6.828157e-17 * -8.398925e-21 = -5.734918e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001100101001000010110111010100;
		b = 32'b01100001010100010110010001000111;
		correct = 32'b01101110100001100100100110111010;
		#400 //86077090.0 * 2.414122e+20 = 2.078006e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010001111100111011001111100111;
		b = 32'b00111000101111101001001011111000;
		correct = 32'b10001011001101010110101101101110;
		#400 //-3.8449513e-28 * 9.087281e-05 = -3.4940153e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001110001111110110100000011001;
		b = 32'b00100110110001110100000011111110;
		correct = 32'b00110101100101001111101010000011;
		#400 //802817600.0 * 1.3826015e-15 = 1.1099768e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100110110000101011001011110110;
		b = 32'b10011001110000000011011001000110;
		correct = 32'b01000001000100100010111101111111;
		#400 //-4.5972017e+23 * -1.9874256e-23 = 9.136596
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111101100011011111101000010100;
		b = 32'b10010000101000111111111010010101;
		correct = 32'b01001110101101011110011011010111;
		#400 //-2.3589953e+37 * -6.468441e-29 = 1525902200.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111100011101010010110011110011;
		b = 32'b11100101100111101110100101111011;
		correct = 32'b11100010100110000011000101011010;
		#400 //0.01496433 * -9.380511e+22 = -1.4037306e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000110010111001110110001000000;
		b = 32'b10010010001001100011001000011011;
		correct = 32'b10011001000011110110110001101111;
		#400 //14139.0625 * -5.2442124e-28 = -7.414825e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111101010101011001001011100110;
		b = 32'b00110110101111110100101010111000;
		correct = 32'b10110100100111111001011011110000;
		#400 //-0.052142046 * 5.700942e-06 = -2.972588e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000111101111001000011101111001;
		b = 32'b10111101101101010000100001000110;
		correct = 32'b01000110000001010101000111100000;
		#400 //-96526.945 * -0.08839469 = 8532.469
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010100101111101001011011100111;
		b = 32'b11010101111110001010111110101111;
		correct = 32'b00101011001110010010010011111011;
		#400 //-1.9244618e-26 * -34179180000000.0 = 6.5776524e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001110010110101010000001001011;
		b = 32'b11100000010111000000011011011110;
		correct = 32'b11101111001110111110011110011110;
		#400 //916984500.0 * -6.3418415e+19 = -5.8153705e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011010111110110011011111001111;
		b = 32'b01111110001101100011101000001101;
		correct = 32'b01011001101100101101001010100101;
		#400 //1.0390133e-22 * 6.055523e+37 = 6291769000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101111010011100011100010011000;
		b = 32'b10111110001101101001110000111100;
		correct = 32'b01101110000100110001101000010111;
		#400 //-6.382233e+28 * -0.17833036 = 1.1381459e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010010010011101101010010010101;
		b = 32'b11001101101111110000010000111100;
		correct = 32'b10100000100110100101010000000111;
		#400 //6.5264166e-28 * -400590720.0 = -2.614422e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100111100111001011111001100101;
		b = 32'b10110101010011100111010000110011;
		correct = 32'b10011101011111001101000010110110;
		#400 //4.3505124e-15 * -7.691007e-07 = -3.3459823e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111111011011011001011101000001;
		b = 32'b11110000110111100100011010000000;
		correct = 32'b01110000110011100100101010011001;
		#400 //-0.9280892 * -5.503272e+29 = 5.1075276e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111000010110011101100000001;
		b = 32'b01111000101111010010000001011101;
		correct = 32'b11110000010011011011100001010011;
		#400 //-8.2987835e-06 * 3.0687516e+34 = -2.5466905e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111101110001000000011001000;
		b = 32'b00010111001000000011110011000000;
		correct = 32'b10001111011001101111100010001011;
		#400 //-2.1994478e-05 * 5.1775466e-25 = -1.1387743e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001101110101110110000011110111;
		b = 32'b11101100100011010000101011111000;
		correct = 32'b11111010111011010101001101000101;
		#400 //451682020.0 * -1.3640827e+27 = -6.1613163e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000010010010101110110100100100;
		b = 32'b11110001111101101110010000101100;
		correct = 32'b01110100110000111011010010111111;
		#400 //-50.731583 * -2.445093e+30 = 1.2404344e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001110100111010010011110010110;
		b = 32'b01010010111000001111110101011110;
		correct = 32'b00100010000010100001111000101101;
		#400 //3.8741608e-30 * 483161740000.0 = 1.8718462e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101100011011001100100100010101;
		b = 32'b10111100011010101110100110011010;
		correct = 32'b01101001010110010100011111011111;
		#400 //-1.1450243e+27 * -0.0143379215 = 1.6417269e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010000000011010101111100100;
		b = 32'b11111011000111101110000100001110;
		correct = 32'b01110101101000001111010000101100;
		#400 //-0.0004946573 * -8.2494756e+35 = 4.0806635e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111100010001001001000111001111;
		b = 32'b10011010101000101000011110001110;
		correct = 32'b11010111011110011001100010110110;
		#400 //4.08259e+36 * -6.722063e-23 = -274434280000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100000110011011101111001101111;
		b = 32'b11000100010100100110101010000101;
		correct = 32'b00100101101010010011011000100000;
		#400 //-3.4875545e-19 * -841.66437 = 2.9353503e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110100000000000100010010100;
		b = 32'b00100000010000101000110000100010;
		correct = 32'b10010111010000101001100100101100;
		#400 //-3.815696e-06 * 1.6478805e-19 = -6.287811e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101100011110011110100011100010;
		b = 32'b11010000101111011010101100100001;
		correct = 32'b11111101101110010010011111111110;
		#400 //1.20848915e+27 * -25456871000.0 = -3.0764354e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011001010111100100101001000101;
		b = 32'b10101101110010000011010111010111;
		correct = 32'b01000111101011011101100011000110;
		#400 //-3910569000000000.0 * -2.2761277e-11 = 89009.55
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000110010101111101100101001110;
		b = 32'b01010010010101011101111000000010;
		correct = 32'b11011001001101000101001011111110;
		#400 //-13814.326 * 229638180000.0 = -3172296700000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111101110000010110100010000010;
		b = 32'b01010110000111010110100011111101;
		correct = 32'b11010100011011011101100011010011;
		#400 //-0.094437614 * 43268560000000.0 = -4086179800000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001110001101000111100101001101;
		b = 32'b11100111011111101110100101101001;
		correct = 32'b11110110001100111011010011100111;
		#400 //756962100.0 * -1.20378674e+24 = -9.11221e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010001011101110100101001001011;
		b = 32'b10010111011101000101011110001010;
		correct = 32'b10101001011011000000011101011111;
		#400 //66381460000.0 * -7.895114e-25 = -5.240892e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110101011100100100001001000011;
		b = 32'b00101110110011000101101111010101;
		correct = 32'b00100100110000010110001110110101;
		#400 //9.024845e-07 * 9.2931586e-11 = 8.386932e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100101011110100001000001110101;
		b = 32'b00101101011000101010111110110000;
		correct = 32'b01010011010111010110111000100100;
		#400 //7.380595e+22 * 1.2885623e-11 = 951035600000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111101001110100100010110000100;
		b = 32'b10100011011011001001110110111010;
		correct = 32'b00100001001011000010101011011010;
		#400 //-0.04547645 * -1.28269855e-17 = 5.833258e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001001011111010100010100101001;
		b = 32'b10101010101010101100110000001100;
		correct = 32'b00110100101010001111100111001100;
		#400 //-1037394.56 * -3.0339652e-13 = 3.147419e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111000110000101100010000010;
		b = 32'b11110011110100010110110010001111;
		correct = 32'b01101011011110010100000110111001;
		#400 //-9.080513e-06 * -3.3184566e+31 = 3.013329e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010110001101011010110100100111;
		b = 32'b11110110001100000010001001101100;
		correct = 32'b11001100111110011111111011110001;
		#400 //1.4675701e-25 * -8.931078e+32 = -131069830.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111110001101011011110001000;
		b = 32'b00001000001001111110101010011001;
		correct = 32'b00010000100000100101011111010100;
		#400 //101743.06 * 5.0530503e-34 = 5.141128e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110001111000111111011100100100;
		b = 32'b11001111101100011000000101111100;
		correct = 32'b11000010000111100001000100101110;
		#400 //6.634666e-09 * -5956106000.0 = -39.516777
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000001010000111110111101100000;
		b = 32'b01010001001001001010000111111000;
		correct = 32'b00010010111111000000001010100010;
		#400 //3.5987587e-38 * 44193250000.0 = 1.5904085e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010111001010010101000001010111;
		b = 32'b11100101111010111101011110110000;
		correct = 32'b00111101100110111111101101100111;
		#400 //-5.470825e-25 * -1.3921686e+23 = 0.076163106
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011010110000011111000111110011;
		b = 32'b01000111000110110001110001101001;
		correct = 32'b00100010011010110000011000001000;
		#400 //8.021382e-23 * 39708.41 = 3.1851632e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011100011111001011101101111001;
		b = 32'b01001110001001101011101001111111;
		correct = 32'b10101011001001001001100110101110;
		#400 //-8.362211e-22 * 699310000.0 = -5.847778e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000100110110101111000011011110;
		b = 32'b01000101011010100111010001100110;
		correct = 32'b11001010110010001000001110110111;
		#400 //-1751.5271 * 3751.275 = -6570459.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000001000011001110010101001111;
		b = 32'b11011001011000011010001111111100;
		correct = 32'b00011010111110000101111110010110;
		#400 //-2.587846e-38 * -3969510800000000.0 = 1.02724823e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101001000111110010101000100100;
		b = 32'b01111001000110110011011011101010;
		correct = 32'b01100010110000010000000101010000;
		#400 //3.5341643e-14 * 5.036999e+34 = 1.7801581e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001010110101000101001001011111;
		b = 32'b10110111110110110100000100010001;
		correct = 32'b11000011001101011101100001101110;
		#400 //6957359.5 * -2.6137133e-05 = -181.84543
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000000010111001010000010101100;
		b = 32'b11010011111011100101111010000010;
		correct = 32'b11010100110011010110111011010011;
		#400 //3.4473066 * -2047575600000.0 = -7058621000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111010000101111011011000110111;
		b = 32'b10101001101010000000010101000110;
		correct = 32'b10100100010001110010010101101000;
		#400 //0.0005787345 * -7.4616135e-14 = -4.318293e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101011100010000011101001010011;
		b = 32'b01000101000100010010011101001000;
		correct = 32'b00110001000110100111101111100000;
		#400 //9.679569e-13 * 2322.455 = 2.2480364e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001010000100011100101011011011;
		b = 32'b11110100100010111110000101001000;
		correct = 32'b00111111000111110101001011100010;
		#400 //-7.019649e-33 * -8.865949e+31 = 0.62235844
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100010011101100110010111111001;
		b = 32'b10100110101011101000100111000000;
		correct = 32'b01001001101001111111110111100101;
		#400 //-1.13631174e+21 * -1.2111013e-15 = 1376188.6
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010101110100010110111110011101;
		b = 32'b11001011000011111000100111100110;
		correct = 32'b00100001011010101101110001010011;
		#400 //-8.459052e-26 * -9406950.0 = 7.957388e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111011000110101111001001001101;
		b = 32'b10110111111010110011100000100101;
		correct = 32'b11110011100011100101111001101000;
		#400 //8.0452816e+35 * -2.8040327e-05 = -2.2559233e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001011001101110001000101001110;
		b = 32'b00111001111110111111010100000101;
		correct = 32'b01000101101101000010110100101111;
		#400 //11997518.0 * 0.00048057004 = 5765.648
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100000010111010000101010101000;
		b = 32'b00100110011010011110000001111101;
		correct = 32'b01000111010010011111000010001000;
		#400 //6.371091e+19 * 8.114235e-16 = 51696.53
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011101000010010111100111100110;
		b = 32'b11110001111100000011001011000011;
		correct = 32'b11001111100000001111110110001010;
		#400 //1.819482e-21 * -2.3788086e+30 = -4328199000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001110000111001011011000011111;
		b = 32'b11011101000000101111011111101110;
		correct = 32'b01101011101000000101100010000010;
		#400 //-657295300.0 * -5.898296e+17 = 3.876922e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010100000101110000100101100;
		b = 32'b01100101011100101010001010101000;
		correct = 32'b11100000011110000001100000001000;
		#400 //-0.0009985319 * 7.1613323e+22 = -7.150819e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110000000001110010110000001;
		b = 32'b10110000011001100100011000111011;
		correct = 32'b00100110111001111110001100011101;
		#400 //-1.9207075e-06 * -8.3773316e-10 = 1.6090404e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111100010110011001101001101111;
		b = 32'b10111100001100000110001100101111;
		correct = 32'b00111001000101011110111001111011;
		#400 //-0.013281449 * -0.010765835 = 0.00014298588
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110111110100100000000001001100;
		b = 32'b00101010000010101010010011100111;
		correct = 32'b00100010011000110111011011011101;
		#400 //2.5034089e-05 * 1.2314074e-13 = 3.0827162e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010000000001011001010011110001;
		b = 32'b00100100110000001111001010000111;
		correct = 32'b10110101010010010101110010000100;
		#400 //-8964523000.0 * 8.3677584e-17 = -7.5012963e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010101011100001011111010010000;
		b = 32'b01011011111100111000101100101111;
		correct = 32'b10110001111001010000011111000110;
		#400 //-4.861794e-26 * 1.3710291e+17 = -6.665661e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000010001001110011111010001001;
		b = 32'b01110011101000010010101000001111;
		correct = 32'b10110110010100101001001110011100;
		#400 //-1.2287169e-37 * 2.5537501e+31 = -3.1378358e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100011100000111100100101010010;
		b = 32'b00101000110011110000111100101111;
		correct = 32'b10001100110101010010111100110101;
		#400 //-1.4288311e-17 * 2.2988201e-14 = -3.2846258e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011111111011000100011010001111;
		b = 32'b01110101110100101111010001011001;
		correct = 32'b01010110010000101011001101100111;
		#400 //1.0006662e-19 * 5.3483315e+32 = 53518946000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011011111011010111110110010110;
		b = 32'b11001110111101101111010000011000;
		correct = 32'b01101011011001010001100100100000;
		#400 //-1.33695305e+17 * -2071596000.0 = 2.7696266e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010110100111001101100010110100;
		b = 32'b01000111000101010011010010111101;
		correct = 32'b00011110001101101101010011100001;
		#400 //2.5339918e-25 * 38196.74 = 9.679022e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011001000110011100010011100101;
		b = 32'b01011011110111110010001011101100;
		correct = 32'b11110101100001100000011101111101;
		#400 //-2705135000000000.0 * 1.2561463e+17 = -3.3980452e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100010011001010100110110110;
		b = 32'b01101010101111100110110100011110;
		correct = 32'b01101111100110000011110100110001;
		#400 //818.65173 * 1.151056e+26 = 9.4231395e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001011010000001010010000000011;
		b = 32'b11101101110011000111011001010010;
		correct = 32'b10111001100110011101101110111100;
		#400 //3.7101244e-32 * -7.909748e+27 = -0.0002934615
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001001000111010111101101111000;
		b = 32'b00110001111010010100100110010101;
		correct = 32'b00111011100011111000001010100100;
		#400 //645047.5 * 6.789558e-09 = 0.0043795872
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011111011011111111011010110110;
		b = 32'b10110010000101110011110011001001;
		correct = 32'b00010010000011011100001110000000;
		#400 //-5.0814293e-20 * -8.803178e-09 = 4.4732727e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100100101110000110110001001101;
		b = 32'b11101110000001110010000100100001;
		correct = 32'b11010011010000101011000111110101;
		#400 //7.998075e-17 * -1.0455132e+28 = -836209300000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111101010001010101101001001011;
		b = 32'b10100110110010101011111001000111;
		correct = 32'b10100100100111000100101111101111;
		#400 //0.048181813 * -1.406814e-15 = -6.778285e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111000100010000000110001101011;
		b = 32'b00110100010101011011101101101001;
		correct = 32'b01101101011000110010101111011100;
		#400 //2.2075132e+34 * 1.990535e-07 = 4.3941325e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001101111010010101000100110110;
		b = 32'b10111000100011001000000111000101;
		correct = 32'b01000111000000000000111010101111;
		#400 //-489301700.0 * -6.699892e-05 = 32782.684
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111111000111101000001011111100;
		b = 32'b10010110011111010010101100001111;
		correct = 32'b10010110000111001100001000011100;
		#400 //0.61918616 * -2.0450764e-25 = -1.266283e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011001001110010000111011000100;
		b = 32'b01101011010011011100011111111001;
		correct = 32'b11000101000101001100000101100001;
		#400 //-9.567258e-24 * 2.4877414e+26 = -2380.0862
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100101110001111110010010000110;
		b = 32'b01010110000100001010110111110110;
		correct = 32'b11111100011000011111000011000010;
		#400 //-1.17995805e+23 * 39769208000000.0 = -4.6925998e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011000101101100000110001110000;
		b = 32'b01011111110111101100111010011001;
		correct = 32'b11111001000111100111000110110100;
		#400 //-1601316300000000.0 * 3.2109876e+19 = -5.1418067e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101001100101110111100101111011;
		b = 32'b00101111100110101001100010110010;
		correct = 32'b00011001101101101111001011011011;
		#400 //6.7268206e-14 * 2.8120933e-10 = 1.8916447e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100010110100000110110000001110;
		b = 32'b01111111001110111001100011111111;
		correct = 32'b11100010100110001011101101111110;
		#400 //-5.649292e-18 * 2.4936004e+38 = -1.4087077e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100000101101100010110010100000;
		b = 32'b11100000100110000011010110111111;
		correct = 32'b01000001110110001010000101111100;
		#400 //-3.086153e-19 * -8.774306e+19 = 27.07885
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111111110101011010110100101001;
		b = 32'b10111011001011001111100011111101;
		correct = 32'b01111111110101011010110100101001;
		#400 //nan * -0.0026393526 = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011100001101101101000101011110;
		b = 32'b11001001011111100011110000010001;
		correct = 32'b10100110001101011000111010100000;
		#400 //6.048935e-22 * -1041345.06 = -6.2990283e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110011110101101101100111111011;
		b = 32'b01000100100010100110000011100001;
		correct = 32'b01111000111010000100010110100000;
		#400 //3.4044577e+31 * 1107.0275 = 3.7688282e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011111000110100010110111101001;
		b = 32'b10101000010011101110111010111011;
		correct = 32'b11000111111110010100000101110010;
		#400 //1.1109792e+19 * -1.14870636e-14 = -127618.89
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101010011011110011100101001011;
		b = 32'b11101110100101110110100010010011;
		correct = 32'b01011001100011010111110010000100;
		#400 //-2.1247342e-13 * -2.342933e+28 = 4978110000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100001101101000110110110001001;
		b = 32'b00000000000100110000110110101011;
		correct = 32'b00100001010101101101110000110100;
		#400 //4.1603835e+20 * 1.749778e-39 = 7.2797457e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001111010010101100100000110100;
		b = 32'b00010101000111111010011110010101;
		correct = 32'b00100100111111001110111000101110;
		#400 //3402118100.0 * 3.2241993e-26 = 1.0969107e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010011010011010100001011011001;
		b = 32'b11000000101000110011000000110110;
		correct = 32'b00010100100000101101100000111000;
		#400 //-2.5907596e-27 * -5.099635 = 1.3211929e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010000110001001001011010100101;
		b = 32'b11000001100100010110011011100010;
		correct = 32'b10010010110111110101000010101010;
		#400 //7.7540473e-29 * -18.175236 = -1.4093164e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100100011001110110111111110010;
		b = 32'b10000000111101101000111010010111;
		correct = 32'b10100101110111101110011001111011;
		#400 //1.7077058e+22 * -2.2642684e-38 = -3.866704e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100010111010110110000011101011;
		b = 32'b00101111111010010000011100000011;
		correct = 32'b00010011010101100100000110101000;
		#400 //6.3799494e-18 * 4.2387435e-10 = 2.7042968e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110100000111110010110111010111;
		b = 32'b10011000101010000010011000111000;
		correct = 32'b01001101010100010001101110110001;
		#400 //-5.044586e+31 * -4.3465573e-24 = 219265810.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001000000100110011001110100110;
		b = 32'b10111000100001011110100010011000;
		correct = 32'b01000001000110011111111100100111;
		#400 //-150734.6 * -6.385258e-05 = 9.624793
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010000101101001010101110100001;
		b = 32'b01111110001010100100001000011111;
		correct = 32'b01001111011100000101000101000110;
		#400 //7.126192e-29 * 5.657802e+37 = 4031858200.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101011111000100111110000101001;
		b = 32'b01011000011100011000011011010010;
		correct = 32'b11000100110101011010111000101001;
		#400 //-1.6092727e-12 * 1062245400000000.0 = -1709.4425
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001110111100110100010010000101;
		b = 32'b00110000100011010001001000110011;
		correct = 32'b11000000000001100000111000001001;
		#400 //-2040677000.0 * 1.0264273e-09 = -2.0946066
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000111101000010100110101010110;
		b = 32'b11111010001100110011111100001101;
		correct = 32'b01000010011000011110000110011011;
		#400 //-2.4270042e-34 * -2.3267499e+35 = 56.470318
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010101100000101000101110100110;
		b = 32'b10110100110100001011000010100010;
		correct = 32'b11001010110101001101011100010011;
		#400 //17942037000000.0 * -3.8871536e-07 = -6974345.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100111100011101001101100001101;
		b = 32'b11001101110100110111011100100100;
		correct = 32'b00110101111010111001100001010100;
		#400 //-3.9581024e-15 * -443475070.0 = 1.7553198e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001010000110010010111111010001;
		b = 32'b00111001110100001100110100101011;
		correct = 32'b00000100011110011110001100111110;
		#400 //7.375675e-33 * 0.00039825714 = 2.9374154e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110101001111011010101000010110;
		b = 32'b11110010001001010000010001001110;
		correct = 32'b01100111111101001000001110100001;
		#400 //-7.0655494e-07 * -3.2684948e+30 = 2.3093711e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101011001001110110010001001111;
		b = 32'b00111001010000100011110000111111;
		correct = 32'b01100100111111100000001011010001;
		#400 //2.023643e+26 * 0.00018523725 = 3.7485408e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100100110000000001010100001101;
		b = 32'b10011111100001010011101111001101;
		correct = 32'b11000100110001111110111110011101;
		#400 //2.8346334e+22 * -5.642662e-20 = -1599.4879
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001001111100010010000001110101;
		b = 32'b10111100100001101101000011111000;
		correct = 32'b01000110111111011111011110100010;
		#400 //-1975310.6 * -0.016457066 = 32507.816
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110100101100101010111010100110;
		b = 32'b11001000111100010011110100000111;
		correct = 32'b10111110001010000110000100000011;
		#400 //3.3282157e-07 * -494056.22 = -0.16443257
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110100111010001000100000001000;
		b = 32'b10101010011111000001001010100111;
		correct = 32'b01011111111001001111011011011001;
		#400 //-1.4738427e+32 * -2.2388568e-13 = 3.2997226e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000001110100100000011111010100;
		b = 32'b11111100011111100010101111111000;
		correct = 32'b00111110110100001000011111010111;
		#400 //-7.715305e-38 * -5.2789408e+36 = 0.40728638
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000011011100111001110111011010;
		b = 32'b01010001001010001011011101001101;
		correct = 32'b01010101001000001000111000000110;
		#400 //243.61661 * 45289360000.0 = 11033240000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110000010001111101000011010;
		b = 32'b11011000001101000100101110101010;
		correct = 32'b11010110110000001111000010101101;
		#400 //0.13376656 * -792948300000000.0 = -106069960000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111001110010010111100011111110;
		b = 32'b11000110000011001000101111010000;
		correct = 32'b01000000010111010011100001100111;
		#400 //-0.00038427854 * -8994.953 = 3.4565675
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110011000000101011110000110000;
		b = 32'b01000000111000000100111001010110;
		correct = 32'b00110100011001010001100101010111;
		#400 //3.043914e-08 * 7.0095625 = 2.1336506e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100000100101101000001000010110;
		b = 32'b10001111000011011001100100000010;
		correct = 32'b00110000001001100111111100110110;
		#400 //-8.676204e+19 * -6.981305e-30 = 6.0571226e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101101100001000001111110010111;
		b = 32'b01000001100110100000100000101110;
		correct = 32'b00101111100111101111111001110011;
		#400 //1.5020691e-11 * 19.253994 = 2.892083e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110010110011011110010001000001;
		b = 32'b10010001110010001100000100111111;
		correct = 32'b01000101001000010111010110111111;
		#400 //-8.156207e+30 * -3.1673533e-28 = 2583.3591
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100110111000110001110010111100;
		b = 32'b11010100100001101000000100010101;
		correct = 32'b11111011111011101010011100011101;
		#400 //5.3625362e+23 * -4621530000000.0 = -2.4783122e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001000101010011101001011110100;
		b = 32'b00001001011001000101101100011100;
		correct = 32'b10010010100101110111110001010010;
		#400 //-347799.62 * 2.7487341e-33 = -9.560087e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110000110100100010001101000100;
		b = 32'b00000011001000000010011111100011;
		correct = 32'b00110100100000110111011011001000;
		#400 //5.202759e+29 * 4.706556e-37 = 2.4487076e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110011100101001011000011101101;
		b = 32'b01011011010010111001110100011110;
		correct = 32'b11001111011011001000011100011100;
		#400 //-6.92397e-08 * 5.7312172e+16 = -3968277500.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101100100111011101000111010000;
		b = 32'b11001011001110101011001100001000;
		correct = 32'b00111000011001100011000110100000;
		#400 //-4.4855022e-12 * -12235528.0 = 5.488249e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011111100101110101011011000110;
		b = 32'b00111000110101101001001111110010;
		correct = 32'b00011000111111011011001111111111;
		#400 //6.409454e-20 * 0.00010231872 = 6.5580717e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010101000010000011001101010001;
		b = 32'b01100101000011000110100001011010;
		correct = 32'b11111010100101010110011100101010;
		#400 //-9359624000000.0 * 4.1441016e+22 = -3.8787232e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111110001100001010010101001;
		b = 32'b00011101100101001100100110101010;
		correct = 32'b00100101111001100011111111110111;
		#400 //101417.32 * 3.938379e-21 = 3.9941984e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100110101000101101101010110;
		b = 32'b01101100010100010001111101011100;
		correct = 32'b01110001101011010111100010010101;
		#400 //1698.8542 * 1.01125435e+27 = 1.7179738e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111101000000010101101011010111;
		b = 32'b00100000101101011100100101110000;
		correct = 32'b01011110001101111011011000000110;
		#400 //1.074638e+37 * 3.0795893e-19 = 3.3094437e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110111000110110110100111010101;
		b = 32'b01101000100011010100010111100001;
		correct = 32'b01100000001010111000011101101101;
		#400 //9.263361e-06 * 5.3371417e+24 = 4.943987e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101011101111100101101110010101;
		b = 32'b00110100100111000111001011001100;
		correct = 32'b01100000111010001010101001010111;
		#400 //4.6025678e+26 * 2.914079e-07 = 1.3412247e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010001001101100110000101000100;
		b = 32'b01111110000011101011101100010110;
		correct = 32'b11001111110010110101111001111001;
		#400 //-1.4387241e-28 * 4.7430445e+37 = -6823932400.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011010000000100110110101110001;
		b = 32'b11100000010111111110111011010111;
		correct = 32'b00111010111001000010111000001001;
		#400 //-2.6971776e-23 * -6.4544284e+19 = 0.0017408739
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001011001110110010011101101010;
		b = 32'b11100001110000111111100001110101;
		correct = 32'b10101101100011110100010010101001;
		#400 //3.6044542e-32 * -4.518773e+20 = -1.6287709e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011101010000110100110101100110;
		b = 32'b10000100000001000011010111000010;
		correct = 32'b10100001110010011011100111010111;
		#400 //8.7956354e+17 * -1.554121e-36 = -1.3669481e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001110111000110111011110010101;
		b = 32'b11110110101101001110000011100110;
		correct = 32'b11000110001000001011011111101010;
		#400 //5.6074974e-30 * -1.834326e+33 = -10285.979
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110100010111011011011010100000;
		b = 32'b10011110010101110110001000010110;
		correct = 32'b01010011001110101000100101010011;
		#400 //-7.0263774e+31 * -1.1402289e-20 = 801167840000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101010010100011011100010010111;
		b = 32'b01111000111110110011010010111000;
		correct = 32'b01100011110011011100101100101100;
		#400 //1.8626971e-13 * 4.0760493e+34 = 7.592445e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100111001110011110000011110101;
		b = 32'b00100011000000010010011110011010;
		correct = 32'b11001010101110111000111000111001;
		#400 //-8.777875e+23 * 7.00149e-18 = -6145820.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111111001000001010111010010010;
		b = 32'b10110100001110011011000000111100;
		correct = 32'b11110011111010010001100110001010;
		#400 //2.135829e+38 * -1.7293581e-07 = -3.6936132e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111100011110000011101000000101;
		b = 32'b00001010010101011000010011111011;
		correct = 32'b00000111010011110000100100110111;
		#400 //0.015150552 * 1.0280588e-32 = 1.5575657e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101011100111111110101110010110;
		b = 32'b10110001101101011011000000111010;
		correct = 32'b10011101111000101111111101001111;
		#400 //1.1363018e-12 * -5.287828e-09 = -6.0085685e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001111110010010000110011011111;
		b = 32'b00101001100011111101111111111110;
		correct = 32'b10111001111000011111110000110101;
		#400 //-6746128000.0 * 6.389332e-14 = -0.00043103253
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011000111011011001001111010100;
		b = 32'b00100010110110011100100101111010;
		correct = 32'b10111100010010100001110101001001;
		#400 //-2089753400000000.0 * 5.903129e-18 = -0.012336084
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101000101000011100100100111111;
		b = 32'b00000110000000000111111100010111;
		correct = 32'b00101111001000100110100111100010;
		#400 //6.1121067e+24 * 2.4167495e-35 = 1.4771431e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000010000011001111110111100000;
		b = 32'b11100010000011011001101011010100;
		correct = 32'b10100100100110111111101000110100;
		#400 //1.0358434e-37 * -6.5303686e+20 = -6.7644395e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110010010111011001100110010001;
		b = 32'b10000110011010010111100110100010;
		correct = 32'b00111001010010100001101000001111;
		#400 //-4.3892376e+30 * -4.391179e-35 = 0.00019273929
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110110110000011101100101101000;
		b = 32'b10101111001001000111100100100011;
		correct = 32'b10100110011110010001011000000010;
		#400 //5.7771576e-06 * -1.495875e-10 = -8.6419055e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100110111100011010100101101101;
		b = 32'b00001010110110000000010000000100;
		correct = 32'b00110010010010111110101010111110;
		#400 //5.7060784e+23 * 2.0801554e-32 = 1.1869529e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011100011101001100001101010101;
		b = 32'b01010101001011001100010101101000;
		correct = 32'b11110010001001010010111111111011;
		#400 //-2.7557866e+17 * 11872741000000.0 = -3.271874e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101011000110100000100011101001;
		b = 32'b11111010111101111101111011011101;
		correct = 32'b01100110100101010010010010110010;
		#400 //-5.4724156e-13 * -6.4350876e+35 = 3.5215476e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011001001001000000000010001110;
		b = 32'b11111100111010001000111001000111;
		correct = 32'b01010110100101001111101110100110;
		#400 //-8.478713e-24 * -9.659989e+36 = 81904270000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110010101110110110101011111000;
		b = 32'b10010010010101111100110011010010;
		correct = 32'b11000101100111011111110011001001;
		#400 //7.424386e+30 * -6.80945e-28 = -5055.598
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101001101001010000111011100101;
		b = 32'b00001100000001111011011011001101;
		correct = 32'b10110110001011110000000101101111;
		#400 //-2.4942887e+25 * 1.0455031e-31 = -2.6077867e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110110101111100100110111001110;
		b = 32'b10110110110111110001000010000110;
		correct = 32'b10101110001001011101001000001111;
		#400 //5.671499e-06 * -6.6478415e-06 = -3.7703226e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101001101000101100010000000101;
		b = 32'b00000000100011111100011111110101;
		correct = 32'b00101010101101101101010101000010;
		#400 //2.4596457e+25 * 1.3204207e-38 = 3.2477672e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010111001010110110110111000011;
		b = 32'b00001111011010101101100000000010;
		correct = 32'b10100111000111010100001011111010;
		#400 //-188487910000000.0 * 1.1578692e-29 = -2.1824435e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100100111010011001001010010110;
		b = 32'b10110110001101011011001010000110;
		correct = 32'b00011011101001011100011110000110;
		#400 //-1.0129597e-16 * -2.7075016e-06 = 2.74259e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010111111111110100000101100111;
		b = 32'b10101110111011001101000000101100;
		correct = 32'b11000111011011000001111111011100;
		#400 //561312730000000.0 * -1.0769016e-10 = -60447.86
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101100000001111111001111110011;
		b = 32'b00100110100000000100100101010101;
		correct = 32'b10010011000010000100000111010110;
		#400 //-1.9320073e-12 * 8.901661e-16 = -1.7198073e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111111100010110010100101000;
		b = 32'b00100000111110101100101101010010;
		correct = 32'b00101001011011000111110010000010;
		#400 //123594.31 * 4.2486193e-19 = 5.251052e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110100001101100111110100001001;
		b = 32'b11101001010100100101001110001111;
		correct = 32'b11011110000101011110111000100010;
		#400 //1.6995558e-07 * -1.5891814e+25 = -2.7009025e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000101010000111010100000001110;
		b = 32'b11011000000111101100011100010001;
		correct = 32'b01011101111100101011001110111011;
		#400 //-3130.5034 * -698311300000000.0 = 2.1860659e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100000100010000111110011110010;
		b = 32'b01101000110111100001011000001000;
		correct = 32'b01001001111011001101000000110010;
		#400 //2.3121978e-19 * 8.390174e+24 = 1939974.2
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011110110000110101100101111100;
		b = 32'b10010001001100101100011000001100;
		correct = 32'b10110000100010000110101101011001;
		#400 //7.038209e+18 * -1.4102752e-28 = -9.925812e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101100010000010000011000111111;
		b = 32'b11100111110100001101110000100000;
		correct = 32'b11010100100111010111101100001101;
		#400 //2.7430417e-12 * -1.9726256e+24 = -5410994500000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111110100000011010001011111;
		b = 32'b10010110100011101010011111110001;
		correct = 32'b10011110111010000000101101000110;
		#400 //106600.74 * -2.3047323e-25 = -2.4568618e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111000011000011100011010011011;
		b = 32'b00100100100101011110011101110100;
		correct = 32'b10011101100001000011010010111001;
		#400 //-5.3829146e-05 * 6.5010546e-17 = -3.4994623e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011001001101100001111111101011;
		b = 32'b00111110100010010011000100111000;
		correct = 32'b01011000010000110011010000110001;
		#400 //3203971200000000.0 * 0.26795363 = 858515700000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010010100001110111001100101001;
		b = 32'b01100110011111001101100111100101;
		correct = 32'b11111001100001011100100010100110;
		#400 //-290876330000.0 * 2.9851395e+23 = -8.683064e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111011101101011011100111100001;
		b = 32'b10100110111111110110100111011101;
		correct = 32'b11100011001101010100111101001101;
		#400 //1.8871516e+36 * -1.7722874e-15 = -3.344575e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111110100101110000001100101001;
		b = 32'b00001001111100011101001100111010;
		correct = 32'b01001001000011101010011010010011;
		#400 //1.0036492e+38 * 5.8217276e-33 = 584297.2
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111010111010110111111001100000;
		b = 32'b11001110010000001111110000101110;
		correct = 32'b11001001101100011000011011000011;
		#400 //0.001796674 * -809438100.0 = -1454296.4
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111001010010111010001100010111;
		b = 32'b10101001101110111111110011010101;
		correct = 32'b11100011100101011000100101000000;
		#400 //6.6084007e+34 * -8.3483276e-14 = -5.5169095e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001011001111100010000110101110;
		b = 32'b00111100110110001101000100110000;
		correct = 32'b10001000101000010000011111001000;
		#400 //-3.6618007e-32 * 0.026466936 = -9.691664e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100001001010110001010110011111;
		b = 32'b10110001110011011010110000101100;
		correct = 32'b00010011100010010111001101100000;
		#400 //-5.796567e-19 * -5.985859e-09 = 3.469743e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011110000011111110110001000011;
		b = 32'b11111001010001000001110100000110;
		correct = 32'b01010111110111001000001001101001;
		#400 //-7.619215e-21 * -6.364243e+34 = 484905330000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001010101101111010101001111110;
		b = 32'b00010000001011001001110001000000;
		correct = 32'b00011011011101111010110101001101;
		#400 //6018367.0 * 3.404139e-29 = 2.0487358e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010101111100101101000100010011;
		b = 32'b01011010001000011111110000100111;
		correct = 32'b11110000100110011010010010101000;
		#400 //-33372473000000.0 * 1.1398679e+16 = -3.804021e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101110111111011001101100111001;
		b = 32'b01100111111010100001110000100010;
		correct = 32'b01010111011001111110101111000001;
		#400 //1.1532681e-10 * 2.2111054e+24 = 254999740000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011110100111101011110101001110;
		b = 32'b10111101011111011100010110001110;
		correct = 32'b01011100100111010101101110010110;
		#400 //-5.719192e+18 * -0.06195598 = 3.5433817e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010101110111110010111001101011;
		b = 32'b11101001111111100111011011101001;
		correct = 32'b11000000010111011101011110111001;
		#400 //9.014222e-26 * -3.8453587e+25 = -3.4662917
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010000110010111101101001111000;
		b = 32'b00101000100010001100111110101011;
		correct = 32'b10111001110110011110001011011011;
		#400 //-27360740000.0 * 1.5189095e-14 = -0.00041558486
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100000010111110010011010100110;
		b = 32'b00110101000000010100111110100111;
		correct = 32'b11010101111000010110111111010000;
		#400 //-6.431889e+19 * 4.8172154e-07 = -30983793000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111111010100100111100100000100;
		b = 32'b01100000001100001001110001010110;
		correct = 32'b01100000000100010011001110111011;
		#400 //0.82215905 * 5.0904565e+19 = 4.185165e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111100000011100011111100110111;
		b = 32'b01000001010110101110010110100001;
		correct = 32'b10111101111100110100001011011010;
		#400 //-0.008682064 * 13.681062 = -0.11877985
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010110111010100101000000010100;
		b = 32'b01011000011011000010110000011001;
		correct = 32'b00101111110110000010101000101111;
		#400 //3.7855275e-25 * 1038696600000000.0 = 3.9320144e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001010110001100011010111000111;
		b = 32'b00101001010001100101110100000111;
		correct = 32'b00110100100110011001010110011111;
		#400 //6494947.5 * 4.404552e-14 = 2.8607334e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011010111100001011100010001100;
		b = 32'b11010000111110110011101100110000;
		correct = 32'b00101100011011000011110010011001;
		#400 //-9.9559825e-23 * -33719680000.0 = 3.3571256e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010101111110100110010100110101;
		b = 32'b11010101111001000100011110010101;
		correct = 32'b01101100010111110100100000100111;
		#400 //-34414073000000.0 * -31374512000000.0 = 1.07972475e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100100010110010000001111101110;
		b = 32'b10011011001110011011000101001110;
		correct = 32'b01000000000111010110101000100101;
		#400 //-1.6012907e+22 * -1.5360132e-22 = 2.4596035
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001100000000010001000110011110;
		b = 32'b10111001010011001100110111111111;
		correct = 32'b10000101110011101000001111001011;
		#400 //9.9431e-32 * -0.00019531696 = -1.942056e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010010111100000111011100010;
		b = 32'b11001001001111010100011101111011;
		correct = 32'b01000100001001000010111011111110;
		#400 //-0.00084708456 * -775287.7 = 656.73425
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011010110010011100110110001000;
		b = 32'b01011100100001001101110100000011;
		correct = 32'b10110111110100010111100001100110;
		#400 //-8.3463705e-23 * 2.991816e+17 = -2.4970806e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000011011111010011111101010111;
		b = 32'b10100000110001010100100100110000;
		correct = 32'b10100100110000110010101000100100;
		#400 //253.24742 * -3.342153e-19 = -8.463916e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001111101100111001101000010011;
		b = 32'b00000010111100111011001001010101;
		correct = 32'b00010011001010101111100001011101;
		#400 //6026438000.0 * 3.5807998e-37 = 2.157947e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000100010110101110011100010;
		b = 32'b11100000100111010011010110001111;
		correct = 32'b01010001101010110010101000111101;
		#400 //-1.013998e-09 * -9.062494e+19 = 91893510000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010000100010011110000011110001;
		b = 32'b00110110100000110011111111000101;
		correct = 32'b10000111100011010110000011101000;
		#400 //-5.438355e-29 * 3.911528e-06 = -2.1272278e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100010111110111000010001101100;
		b = 32'b01110111110011110001000011100111;
		correct = 32'b01011011010010110111000010101111;
		#400 //6.8173893e-18 * 8.399596e+33 = 5.7263317e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110100100110001111111101111000;
		b = 32'b00101110001000011111110100000110;
		correct = 32'b01100011010000011001111111000101;
		#400 //9.697396e+31 * 3.683189e-11 = 3.5717342e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100000001111100010001000101101;
		b = 32'b11001010000111100110111011001010;
		correct = 32'b10101010111010110101011011000001;
		#400 //1.6104934e-19 * -2595762.5 = -4.1804583e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001001000110110111011011010001;
		b = 32'b01001010001001010101110100100001;
		correct = 32'b01010011110010001101100001000110;
		#400 //636781.06 * 2709320.2 = 1725243900000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000000101110100100100100101100;
		b = 32'b00011110100110100101010100100110;
		correct = 32'b10011111111000001001101111110101;
		#400 //-5.821432 * 1.63406e-20 = -9.51257e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010100110110000100101100111000;
		b = 32'b00101001111000010110101101101010;
		correct = 32'b10111111001111100111010011011101;
		#400 //-7431799000000.0 * 1.00106406e-13 = -0.7439707
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011100110110010111001010110101;
		b = 32'b01110100101010001110000101011010;
		correct = 32'b01010010000011110111001010110001;
		#400 //1.4389507e-21 * 1.0704059e+32 = 154026130000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100110011111001110001100100011;
		b = 32'b11111101111100000001111111011011;
		correct = 32'b11100100111011010011010001101001;
		#400 //8.773789e-16 * -3.9897515e+37 = -3.500524e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111001111101110101110110101;
		b = 32'b11010111000010111111110010011111;
		correct = 32'b01001110110100001100110011000100;
		#400 //-1.1379762e-05 * -153917120000000.0 = 1751540200.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000001000010010001001001101110;
		b = 32'b10111010010110111110101001111101;
		correct = 32'b10111011111010111000000010100100;
		#400 //8.566999 * -0.00083891285 = -0.007186966
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011101000111010001100100110010;
		b = 32'b00100011000011100111010011001100;
		correct = 32'b10000000101011101101011101001101;
		#400 //-2.0791803e-21 * 7.722568e-18 = -1.6056612e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111101011100001010011011010111;
		b = 32'b11000000010111110011001100101010;
		correct = 32'b10111110010100011101000101101110;
		#400 //0.05875286 * -3.4874978 = -0.20490047
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111101100111001000010000100100;
		b = 32'b00111001111110110101001011011010;
		correct = 32'b11111000000110011010100000110111;
		#400 //-2.600571e+37 * 0.0004793618 = -1.2466144e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110101100101000001001000000010;
		b = 32'b01101111000000100010110111101001;
		correct = 32'b11100101000101101001011101100110;
		#400 //-1.10321e-06 * 4.0288553e+28 = -4.4446736e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000100111100011011101011011000;
		b = 32'b01001101001010011000100001011000;
		correct = 32'b11010010101000000001010100010111;
		#400 //-1933.8389 * 177767800.0 = -343774300000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000011001101110011110111111000;
		b = 32'b11111010111011001111011111001111;
		correct = 32'b01111110101010011001111010000010;
		#400 //-183.24207 * -6.152041e+35 = 1.1273128e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011101101111100110110001011111;
		b = 32'b11000010001010000010110000100100;
		correct = 32'b10100000011110100010111111100111;
		#400 //5.0404634e-21 * -42.043106 = -2.1191673e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011101000000111101000110100001;
		b = 32'b00011010001011111110101110001110;
		correct = 32'b10110111101101010010101100101111;
		#400 //-5.936594e+17 * 3.637943e-23 = -2.159699e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101101111100110110101110001011;
		b = 32'b01001000101010001010000111010011;
		correct = 32'b00110111001000000101100001110010;
		#400 //2.767366e-11 * 345358.6 = 9.557336e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010101101110000000111010111001;
		b = 32'b10111001000101100010100110010100;
		correct = 32'b00001111010101111110110100001010;
		#400 //-7.4340236e-26 * -0.00014320604 = 1.06459705e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011001001110111001110010111100;
		b = 32'b01010011000101010101100111001011;
		correct = 32'b01101100110110101110100000001111;
		#400 //3300509500000000.0 * 641456600000.0 = 2.1171336e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011001010111110000110110001101;
		b = 32'b01100100100100100010000100001111;
		correct = 32'b10111110011111101010010100010000;
		#400 //-1.1531566e-23 * 2.1564854e+22 = -0.24867654
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010100111110000011000101000101;
		b = 32'b00101110101011101111101101010010;
		correct = 32'b00000100001010011010010100100101;
		#400 //2.5061034e-26 * 7.9572474e-11 = 1.9941685e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011011101000001011010101001011;
		b = 32'b10111111000110110000010110011100;
		correct = 32'b00011011010000101010001010010100;
		#400 //-2.6586937e-22 * -0.60555434 = 1.6099836e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001110111010111011010101001010;
		b = 32'b11011011110101010000000111111111;
		correct = 32'b11101011010001000001111110101101;
		#400 //1977263400.0 * -1.1991273e+17 = -2.3709905e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011001011001001010111000000011;
		b = 32'b11011111110110110111111000111100;
		correct = 32'b10111001110001000001000110100000;
		#400 //1.1822465e-23 * -3.163229e+19 = -0.00037397165
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111111001011110010011001001100;
		b = 32'b11000011111110101011011011011111;
		correct = 32'b01000011101010111000100010000100;
		#400 //-0.6841781 * -501.42868 = 343.06653
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010100010100100111111010010110;
		b = 32'b10110001011000101010010111010101;
		correct = 32'b00000110001110100101110000011011;
		#400 //-1.0627255e-26 * -3.2981593e-09 = 3.505038e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000011011000001011001001111110;
		b = 32'b00011100110110101001001101000011;
		correct = 32'b10100000101111111101100101000001;
		#400 //-224.69724 * 1.4464096e-21 = -3.2500425e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011010100101010011101110100011;
		b = 32'b00111101010110000100110011011111;
		correct = 32'b00011000011111000010111001000010;
		#400 //6.1721304e-23 * 0.052807685 = 3.259359e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010100001001001010001000001111;
		b = 32'b11001101111001100001100101101101;
		correct = 32'b00100010100100111111100111110011;
		#400 //-8.3118445e-27 * -482553250.0 = 4.0109074e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100101011111001101010010001000;
		b = 32'b00001001100100110100010100001110;
		correct = 32'b10101111100100010111001000111101;
		#400 //-7.4622304e+22 * 3.54539e-33 = -2.6456518e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001001011101100011001110100011;
		b = 32'b11100001011010111011011011000110;
		correct = 32'b01101011011000101011000100101110;
		#400 //-1008442.2 * -2.717597e+20 = 2.7405394e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110101000101100000110110110100;
		b = 32'b01010000001001100111110000010100;
		correct = 32'b01000101110000110010101100111010;
		#400 //5.5899295e-07 * 11172598000.0 = 6245.4033
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001110101011101100011010011100;
		b = 32'b00011100011011101010101101010111;
		correct = 32'b00101011101000101111000110011111;
		#400 //1466125800.0 * 7.8969046e-22 = 1.1577856e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100100110101111000011010000011;
		b = 32'b00110000011101011011010110000111;
		correct = 32'b10010101110011101101110010001111;
		#400 //-9.346926e-17 * 8.9388447e-10 = -8.355072e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110110101101001101001110000000;
		b = 32'b11100000010010101001000001100111;
		correct = 32'b11010111100011110001010011100011;
		#400 //5.38904e-06 * -5.838512e+19 = -314639740000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000101000100011011101001110111;
		b = 32'b01010110011101111110111110111001;
		correct = 32'b01011100000011010010001101011111;
		#400 //2331.654 * 68152243000000.0 = 1.5890745e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100110101100101001000111010001;
		b = 32'b10010001001111111101011111000100;
		correct = 32'b10111000100001011101000101001100;
		#400 //4.2163554e+23 * -1.5133731e-28 = -6.380919e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000001011111111111010110011011;
		b = 32'b11100100101100010111111000101101;
		correct = 32'b10100110101100010111011011111000;
		#400 //4.7012316e-38 * -2.6193325e+22 = -1.2314089e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010111110011111111001111010000;
		b = 32'b00001110001110010111101110100101;
		correct = 32'b10100110100101101010101110100001;
		#400 //-457292150000000.0 * 2.2862543e-30 = -1.0454861e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010001100110101101001100100011;
		b = 32'b11010010001110000011010110011011;
		correct = 32'b01100100010111101101000001011001;
		#400 //-83120910000.0 * -197793330000.0 = 1.6440761e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010011100011000111101100110010;
		b = 32'b00111110000100001001111110101000;
		correct = 32'b11010010000111101011100111010010;
		#400 //-1206724600000.0 * 0.14123404 = -170430600000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001101110011010100111100110000;
		b = 32'b00111011100111101000101110010101;
		correct = 32'b11001001111111100100110110100010;
		#400 //-430564860.0 * 0.004838417 = -2083252.2
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001110011001101000001111101101;
		b = 32'b11010110110010000010011101010001;
		correct = 32'b10100101101101000011101001111000;
		#400 //2.8413209e-30 * -110035590000000.0 = -3.1264643e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010000110111110010101110100000;
		b = 32'b11000010111010100000001011011110;
		correct = 32'b01010100010011000000000001100000;
		#400 //-29953425000.0 * -117.0056 = 3504718500000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101011000100001001001000001010;
		b = 32'b00000000100010101010000010010110;
		correct = 32'b10101100000111001001001011010011;
		#400 //-1.7477497e+26 * 1.2730906e-38 = -2.2250437e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010111110101100000110001101110;
		b = 32'b10111100010010001100110000110101;
		correct = 32'b11010100101001111110010001110100;
		#400 //470697750000000.0 * -0.012255718 = -5768739000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010111111011011000010010011111;
		b = 32'b00101101101011110000001101000100;
		correct = 32'b01000110001000100110000010110000;
		#400 //522307720000000.0 * 1.9896647e-11 = 10392.172
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110110000101101000111101001100;
		b = 32'b10111100010000110010000110010001;
		correct = 32'b01110010111001011000010111001001;
		#400 //-7.6342865e+32 * -0.011909858 = 9.092327e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111011000101110010010111010101;
		b = 32'b00011000110101101110000111101100;
		correct = 32'b00010100011111011011111000000111;
		#400 //0.002306332 * 5.5545826e-24 = 1.2810712e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111010011110011010100000111001;
		b = 32'b01010001000101101101011110111001;
		correct = 32'b01001100000100110001101011110010;
		#400 //0.00095236633 * 40491520000.0 = 38562760.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100001100001001011111100110110;
		b = 32'b01001011100011001000110000101010;
		correct = 32'b00101101100100011100001010000000;
		#400 //8.995281e-19 * 18421844.0 = 1.6570967e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100010010101100000010011000010;
		b = 32'b11100101100110010110001100101101;
		correct = 32'b11001000100000000011101111000001;
		#400 //2.9004927e-18 * -9.054394e+22 = -262622.03
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000010100101110000101110011101;
		b = 32'b01110100011110100010011111001110;
		correct = 32'b10110111100100111001100011010100;
		#400 //-2.2194122e-37 * 7.927744e+31 = -1.7594932e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000111101011001000000001111100;
		b = 32'b11010100111000101111111110100110;
		correct = 32'b01011101000110001111010110110001;
		#400 //-88320.97 * -7799613400000.0 = 6.888694e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000111001110110101110110101001;
		b = 32'b01101000100111011101001010001010;
		correct = 32'b00110000011001110000010100010001;
		#400 //1.4095841e-34 * 5.9623624e+24 = 8.404451e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110011100111000111100100001110;
		b = 32'b00111010001100111101001110011000;
		correct = 32'b10101110010110111101001111110011;
		#400 //-7.286336e-08 * 0.0006859838 = -4.9983084e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000010111101011010110001000011;
		b = 32'b11001010011010100001010001101101;
		correct = 32'b00001101111000001010001100001111;
		#400 //-3.6098388e-37 * -3835163.2 = 1.3844321e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000111001110010001110110011000;
		b = 32'b01000000110111001011010011110000;
		correct = 32'b10001000100111111001100001000101;
		#400 //-1.392655e-34 * 6.897087 = -9.605263e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011011011010001110000111001111;
		b = 32'b01001001111011110001010011001001;
		correct = 32'b10100101110110010111110110111001;
		#400 //-1.9263553e-22 * 1958553.1 = -3.7728692e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100110010110101110000001000001;
		b = 32'b01101101010010101000111100001000;
		correct = 32'b01010100001011010010111100111101;
		#400 //7.5937864e-16 * 3.9180554e+27 = 2975287500000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000111000111101011100101000000;
		b = 32'b11001001100001100000111001001100;
		correct = 32'b10010001001001100011101110101010;
		#400 //1.1941039e-34 * -1098185.5 = -1.3113476e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100011100011101111101111100110;
		b = 32'b01011000001100110011011010011000;
		correct = 32'b11111100010010000011000101000000;
		#400 //-5.2751777e+21 * 788188240000000.0 = -4.157833e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001000010110110001011100010111;
		b = 32'b11101000010100000010101110101100;
		correct = 32'b00110001001100100010100000100011;
		#400 //-6.5930057e-34 * -3.9322313e+24 = 2.5925224e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100100000111111011110000100010;
		b = 32'b00110010110000101110110110111111;
		correct = 32'b10010111011100110100000111010100;
		#400 //-3.4636984e-17 * 2.2692687e-08 = -7.860062e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111000010100111000000101100000;
		b = 32'b00100000101000110001110101001100;
		correct = 32'b10011001100001101100001110010101;
		#400 //-5.042681e-05 * 2.763266e-19 = -1.393427e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110000110001111111101011111011;
		b = 32'b11000010100110010000101010101011;
		correct = 32'b01110011111011110001101010101011;
		#400 //-4.9512747e+29 * -76.520836 = 3.7887568e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101001000101010000001101110110;
		b = 32'b11100101010001001110010010001111;
		correct = 32'b11001110111001010011011101100001;
		#400 //3.3087648e-14 * -5.81125e+22 = -1922805900.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111011101110110101110011010100;
		b = 32'b00010111001111101011100111010101;
		correct = 32'b01010011100010111001011011100111;
		#400 //1.9456846e+36 * 6.1626864e-25 = 1199064400000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001011010101101010101010111001;
		b = 32'b01100011101010100001000011101000;
		correct = 32'b00101111100011101001101110001100;
		#400 //4.1343338e-32 * 6.2743294e+21 = 2.5940172e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011101001000010011101000001000;
		b = 32'b11111101010111101100010001000001;
		correct = 32'b11011011000011000100101111101100;
		#400 //2.1338174e-21 * -1.8506726e+37 = -3.9489974e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001011010111000000100011101110;
		b = 32'b11000110001101000001001011011101;
		correct = 32'b00010010000110101100011001111110;
		#400 //-4.2377177e-32 * -11524.716 = 4.883849e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001110101111110110100110010101;
		b = 32'b11100111001011010100101011111110;
		correct = 32'b00110110100000011001001001101100;
		#400 //-4.7186807e-30 * -8.1835276e+23 = 3.8615453e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000110101111101011011100000101;
		b = 32'b00000111011100100010001010011010;
		correct = 32'b00001110101101000110001011001010;
		#400 //24411.51 * 1.8216225e-34 = 4.4468556e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100010010110010100001011111011;
		b = 32'b10100000011110101101100011000100;
		correct = 32'b01000011010101001110001101100000;
		#400 //-1.0019425e+21 * -2.1247545e-19 = 212.88818
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001000100111011010111011101000;
		b = 32'b10010001010010100000000010111101;
		correct = 32'b00011010011110001101100011101111;
		#400 //-322935.25 * -1.5935218e-28 = 5.1460436e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011000100111100100011011100010;
		b = 32'b01101010101011001110011110101011;
		correct = 32'b11000011110101011100110110110111;
		#400 //-4.0913616e-24 * 1.0451463e+26 = -427.60715
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011101001101110001010101001110;
		b = 32'b11110110110101100110000001011101;
		correct = 32'b11010100100110010101000010111010;
		#400 //2.4230863e-21 * -2.1740352e+33 = -5267875000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111110000011110111010101010001;
		b = 32'b00100111110110011001010100011000;
		correct = 32'b10100110011100111101101111111101;
		#400 //-0.14009596 * 6.0391247e-15 = -8.46057e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010110100000110111101111010;
		b = 32'b01100100000110111110010111111001;
		correct = 32'b11011111011111011101110101111011;
		#400 //-0.0015902363 * 1.1503266e+22 = -1.8292913e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011110010011100110001000100110;
		b = 32'b00110101010100111010001010010001;
		correct = 32'b01010100001010101001110111110100;
		#400 //3.7178727e+18 * 7.884019e-07 = 2931177800000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001111010001000111001110010001;
		b = 32'b11001111010110011000001001001111;
		correct = 32'b11011111001001101110100111110101;
		#400 //3295908000.0 * -3649195800.0 = -1.2027414e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110010110000001000000101101110;
		b = 32'b10010000001001101010110110101100;
		correct = 32'b10000011011110101010110100001100;
		#400 //2.24106e-08 * -3.287152e-29 = -7.3667045e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110010110110001100101000111101;
		b = 32'b10010011111011000010111010010001;
		correct = 32'b00000111010010000000000111011111;
		#400 //-2.5237677e-08 * -5.9620694e-27 = 1.5046878e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001110111110110111101011000101;
		b = 32'b11001000111010010011000111001001;
		correct = 32'b01011000011001010001001110100101;
		#400 //-2109563500.0 * -477582.28 = 1007490140000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000101100101001110011110000011;
		b = 32'b10110001000000011011101011000010;
		correct = 32'b00110111000101101110101010010100;
		#400 //-4764.939 * -1.887813e-09 = 8.995314e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100110110101011000111111000010;
		b = 32'b00011101011010011101011110010001;
		correct = 32'b00000100110000110001001110101100;
		#400 //1.481881e-15 * 3.0948738e-21 = 4.5862345e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011011000010101010111010100001;
		b = 32'b10110001010010111100011011110001;
		correct = 32'b10001100110111001100100001111111;
		#400 //1.1471518e-22 * -2.9653473e-09 = -3.4017036e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101010000110100110100111011010;
		b = 32'b01111111010100111110010010110100;
		correct = 32'b11101001111111111001111001100011;
		#400 //-1.3714672e-13 * 2.816546e+38 = -3.8628006e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011010111111111000011000010111;
		b = 32'b00100000010000100101011101111010;
		correct = 32'b10111011110000011111101011101110;
		#400 //-3.5961776e+16 * 1.6461383e-19 = -0.0059198057
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100101000111010111101100011011;
		b = 32'b11010000110010011001000011100110;
		correct = 32'b01110110011101111111110110010110;
		#400 //-4.648015e+22 * -27053732000.0 = 1.2574616e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110110111000010100000101001;
		b = 32'b11000100100011011001100110011000;
		correct = 32'b11000011111100111000110001101011;
		#400 //0.4299939 * -1132.7998 = -487.09702
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110001010000111010111000101;
		b = 32'b10100010000001110111100110011100;
		correct = 32'b00011000101100100100110001000010;
		#400 //-2.5102502e-06 * -1.8360291e-18 = 4.6088922e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010100100110001000110000110011;
		b = 32'b11010000110010011000110000110001;
		correct = 32'b01100101111100000011001100111100;
		#400 //-5241497500000.0 * -27051264000.0 = 1.4178913e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001000001101111110010011100010;
		b = 32'b11001011111110010010101111000111;
		correct = 32'b11010100101100101111110100010010;
		#400 //188307.53 * -32659342.0 = -6150000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101110001011111010011110110010;
		b = 32'b00010111001110011000110111001101;
		correct = 32'b01000101111111101010001011110111;
		#400 //1.3590652e+28 * 5.99557e-25 = 8148.3706
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010001111010100010010100100010;
		b = 32'b00001110111101100011011101001110;
		correct = 32'b00100001011000010011001001000100;
		#400 //125705670000.0 * 6.069694e-30 = 7.629949e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010110101101100011101100000001;
		b = 32'b01010010100001000000100100011110;
		correct = 32'b00101001101110111111100111010100;
		#400 //2.9440923e-25 * 283544320000.0 = 8.3478065e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110100101010010111111101011111;
		b = 32'b11010101100001100100111000111111;
		correct = 32'b01001010101100011101100011110100;
		#400 //-3.1571378e-07 * -18458828000000.0 = 5827706.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110100111000111100000011110100;
		b = 32'b11101100011010101110001011110111;
		correct = 32'b01100001110100001111100001001011;
		#400 //-4.2422437e-07 * -1.1358418e+27 = 4.8185177e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001100010010110111100001001000;
		b = 32'b01010110111010100011111101100011;
		correct = 32'b10100011101110100010111001010011;
		#400 //-1.5674747e-31 * 128778980000000.0 = -2.018578e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100010101101101001110111011111;
		b = 32'b11000110111101111000001100011101;
		correct = 32'b11101010001100001000111111011010;
		#400 //1.6843416e+21 * -31681.557 = -5.3362566e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101111000101110011011101110000;
		b = 32'b01001100011101111110100011010011;
		correct = 32'b01111100000100100111000000000100;
		#400 //4.6799256e+28 * 64987980.0 = 3.041389e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010101010010011011010100001101;
		b = 32'b01100110000000000101101100011101;
		correct = 32'b01111011110010100100010010100001;
		#400 //13861215000000.0 * 1.5153591e+23 = 2.1004719e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000011101110011000001010001000;
		b = 32'b00101111010011110110000110111110;
		correct = 32'b00110011100101100100011101100000;
		#400 //371.01978 * 1.8861265e-10 = 6.997902e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100111011111010101101110000001;
		b = 32'b10101110011010010000001001111101;
		correct = 32'b01010110011001101001101010111111;
		#400 //-1.1964467e+24 * -5.2980276e-11 = 63388076000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010110110101011011010010001011;
		b = 32'b00001111110001001000000011010101;
		correct = 32'b00100111001001000000100111000111;
		#400 //117485700000000.0 * 1.9376716e-29 = 2.2764872e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010111110010111101101010111100;
		b = 32'b10100111010110011010101010011011;
		correct = 32'b10111111101011010101010001000100;
		#400 //448280630000000.0 * -3.0207285e-15 = -1.3541341
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000001001010111111100110010011;
		b = 32'b11101110011100101111011111000101;
		correct = 32'b10110000001000110011100001011111;
		#400 //3.15868e-38 * -1.8798727e+28 = -5.937916e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010111101010011010001100001100;
		b = 32'b11111000110101010101111101011100;
		correct = 32'b01010001000011010110001111011001;
		#400 //-1.0962528e-24 * -3.4621667e+34 = 37954097000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111010001111100011101011111110;
		b = 32'b00100110110100110000100011110111;
		correct = 32'b00100001100111001101000101001001;
		#400 //0.00072567153 * 1.4643496e-15 = 1.0626369e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010011011010001000010100011001;
		b = 32'b10110101111101000011010011011010;
		correct = 32'b01001001110111011100111011011101;
		#400 //-998665400000.0 * -1.8194798e-06 = 1817051.6
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001100000110110000111000000010;
		b = 32'b11010101001010100100101011100101;
		correct = 32'b00100001110011100100100101010100;
		#400 //-1.1944981e-31 * -11702415000000.0 = 1.3978513e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110110110011010011111101011101;
		b = 32'b01000001111001110010011100011011;
		correct = 32'b00111001001110010101001110000111;
		#400 //6.1168525e-06 * 28.894094 = 0.00017674091
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111100011010101100001110000000;
		b = 32'b10111111010011100001110100010000;
		correct = 32'b00111100001111010000001111111000;
		#400 //-0.014328837 * -0.80513096 = 0.011536591
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000010100011010100010101110001;
		b = 32'b11000000101100101011010101100110;
		correct = 32'b10000011110001010011110011000110;
		#400 //2.0757945e-37 * -5.5846434 = -1.1592572e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011001011011011110001011111000;
		b = 32'b01001000101000110111110010100011;
		correct = 32'b01100010100101111110101101010101;
		#400 //4184945300000000.0 * 334821.1 = 1.4012079e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101110010010101011110010010000;
		b = 32'b00111100110010000111101110101111;
		correct = 32'b11101011100111101100010101000100;
		#400 //-1.5685983e+28 * 0.02447304 = -3.8388368e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010000100101001010011100001011;
		b = 32'b11100110111001000010111011100010;
		correct = 32'b10111000000001000111111111111111;
		#400 //5.863308e-29 * -5.387822e+23 = -3.1590458e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001100110011110001011010111011;
		b = 32'b01011010101001111010110001110110;
		correct = 32'b10101000000001111010001101010111;
		#400 //-3.190708e-31 * 2.3597972e+16 = -7.529424e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100010101100110101100001011101;
		b = 32'b01011100000110000010001100111011;
		correct = 32'b01111111010101010010101001001011;
		#400 //1.6541672e+21 * 1.7129173e+17 = 2.8334516e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011011000111111000100100100011;
		b = 32'b11001000101110001111011110010111;
		correct = 32'b01100100011001101000100110111001;
		#400 //-4.4905305e+16 * -378812.72 = 1.70107e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001101100001110101000100111100;
		b = 32'b11001100100111001110011110010011;
		correct = 32'b00011010101001011101111111010001;
		#400 //-8.339574e-31 * -82263190.0 = 6.8603995e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101100100100001011100010110110;
		b = 32'b00100111010001000011000100110001;
		correct = 32'b00010100010111011101001001110101;
		#400 //4.113233e-12 * 2.722713e-15 = 1.1199154e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001111000010101111101010011010;
		b = 32'b01100010111110011110001000101101;
		correct = 32'b00110010100001111010100010001001;
		#400 //6.8521894e-30 * 2.3047685e+21 = 1.579271e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101011100111101100011000100110;
		b = 32'b00110101000100100000001101101000;
		correct = 32'b11100001001101010001111000111101;
		#400 //-3.83892e+26 * 5.4394195e-07 = -2.0881497e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110011100100000001111001101000;
		b = 32'b11001010010111001110010010100110;
		correct = 32'b10111110011110001011010110110100;
		#400 //6.7110534e-08 * -3619113.5 = -0.24288064
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100010100100110011001100101101;
		b = 32'b10100000011001000100110110101110;
		correct = 32'b10000011100000110100011000111111;
		#400 //3.9898614e-18 * -1.9338053e-19 = -7.715616e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100101101111111001100110101000;
		b = 32'b00001101010010110011000100010001;
		correct = 32'b10110011100110000001001110010001;
		#400 //-1.1310081e+23 * 6.2613266e-31 = -7.081611e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101000101010011101010011000100;
		b = 32'b10001100000010100010110101001100;
		correct = 32'b10110101001101110101010101111101;
		#400 //6.416038e+24 * -1.0644764e-31 = -6.8297214e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011011000010110111100110101001;
		b = 32'b01000001010100010111101000001001;
		correct = 32'b11011100111001000100000110100000;
		#400 //-3.925879e+16 * 13.092294 = -5.139876e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100111001111010101101100000;
		b = 32'b10000011100001000011101000000101;
		correct = 32'b10001000111011110101000110111110;
		#400 //1853.3555 * -7.771583e-37 = -1.4403507e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100101011110001110111000100010;
		b = 32'b00011000001100010111001110011001;
		correct = 32'b00111110001011001000110100001101;
		#400 //7.347123e+22 * 2.2935076e-24 = 0.16850682
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010101101010010000001011111010;
		b = 32'b10101110000100110100100011111011;
		correct = 32'b11000100010000100111100111001000;
		#400 //23228781000000.0 * -3.348875e-11 = -777.90283
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101011111111010100001001110100;
		b = 32'b01101100111100111001101010110101;
		correct = 32'b01011001011100001111111100100001;
		#400 //1.7995176e-12 * 2.3559965e+27 = 4239657000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110001101011001010100011110001;
		b = 32'b00101110100100101001100101110000;
		correct = 32'b10100000110001011011111110101100;
		#400 //-5.0250653e-09 * 6.666567e-11 = -3.3499936e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010010100110000001010010001001;
		b = 32'b00111010100100100101101101001110;
		correct = 32'b10001101101011011110001111101000;
		#400 //-9.597611e-28 * 0.0011166127 = -1.0716815e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010110000101100110100010000011;
		b = 32'b00000000101100100001000000100101;
		correct = 32'b10010111010100010011110001001111;
		#400 //-41343905000000.0 * 1.635251e-38 = -6.760766e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110011110111001000010000001111;
		b = 32'b00000001011101001111110110110010;
		correct = 32'b00110101110100110000100001100110;
		#400 //3.4942132e+31 * 4.499774e-38 = 1.5723169e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111110111101101100011111111101;
		b = 32'b00001000110000011111101001110101;
		correct = 32'b11001000001110101111111000110110;
		#400 //-1.6401424e+38 * 1.1674647e-33 = -191480.84
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100001101111110001010011001001;
		b = 32'b10011010011110001010100101001111;
		correct = 32'b10111100101110011001101010000010;
		#400 //4.4060323e+20 * -5.1421964e-23 = -0.022656683
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100100000101011110100010011000;
		b = 32'b01001110010111100000111001000001;
		correct = 32'b00110011000000100000100000001101;
		#400 //3.250624e-17 * 931369000.0 = 3.0275306e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110011111110001011110000100;
		b = 32'b11101001011100010101101011010111;
		correct = 32'b01100000011100000111111110101000;
		#400 //-3.801165e-06 * -1.8236256e+25 = 6.931902e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101100001010001011000111000001;
		b = 32'b01110111100011010100100000111000;
		correct = 32'b11100100001110100011001011111100;
		#400 //-2.397291e-12 * 5.731083e+33 = -1.3739073e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110001110100101110100010100110;
		b = 32'b10111000001011010010101000100010;
		correct = 32'b00101010100011101010100111101110;
		#400 //-6.1382535e-09 * -4.1285653e-05 = 2.534218e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000010000000001010100101111111;
		b = 32'b11100011011010001000011111010110;
		correct = 32'b10100101111010011011101111000000;
		#400 //9.452598e-38 * -4.2894326e+21 = -4.0546281e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011011000110001110101000000100;
		b = 32'b01000111100010100111010000001101;
		correct = 32'b11100011001001010110011011110000;
		#400 //-4.30415e+16 * 70888.1 = -3.0511302e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100100011010111100101110001010;
		b = 32'b10001110110010001100110111101001;
		correct = 32'b00110011101110001111010010101100;
		#400 //-1.7398606e+22 * -4.950209e-30 = 8.612673e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011011100011000110100011111110;
		b = 32'b10111000010000011000110010000101;
		correct = 32'b11010100010101000101000001110100;
		#400 //7.904387e+16 * -4.6145655e-05 = -3647531400000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001101101011001000011101011011;
		b = 32'b01000111100000000010100011100010;
		correct = 32'b00010101101011001011111001110110;
		#400 //1.0632904e-30 * 65617.766 = 6.977074e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111001101100010101101010000001;
		b = 32'b01010001101100100101010011111111;
		correct = 32'b01001011111101110001011110100000;
		#400 //0.00033827501 * 95741270000.0 = 32386880.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101000000010000100000010111101;
		b = 32'b00011110000000000101101100001011;
		correct = 32'b10000110100010001010000110100111;
		#400 //-7.5635544e-15 * 6.795091e-21 = -5.139504e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100011001101110011101011110100;
		b = 32'b11011011000000010011011010010101;
		correct = 32'b01111110101110001111011110001100;
		#400 //-3.3800022e+21 * -3.6370286e+16 = 1.2293164e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010000000000110001010010001000;
		b = 32'b11100010000000100111011001010001;
		correct = 32'b00110010100001011001101000000100;
		#400 //-2.585101e-29 * -6.016506e+20 = 1.5553276e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100011000100011111111110000110;
		b = 32'b00111101110100101101010010101111;
		correct = 32'b10100001011100000111100111001111;
		#400 //-7.914575e-18 * 0.102944724 = -8.1476375e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110100111111101111010110110110;
		b = 32'b00101010100010000101010000000010;
		correct = 32'b11100000000001111100011000110011;
		#400 //-1.6159998e+32 * 2.4216745e-13 = -3.9134253e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111111111111101101000100111111;
		b = 32'b10111001000010100110001011001110;
		correct = 32'b10111001100010011011111100100101;
		#400 //1.9907607 * -0.00013197513 = -0.0002627309
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111101101111100111110011110111;
		b = 32'b10001010001100011101000110000111;
		correct = 32'b10001000100001000101000001001111;
		#400 //0.09301179 * -8.561648e-33 = -7.9633415e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111011000111011000010001101010;
		b = 32'b10110001111010111111010111001111;
		correct = 32'b10101101100100010010111111001100;
		#400 //0.0024035224 * -6.8673454e-09 = -1.6505818e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001110101110010001001111000101;
		b = 32'b11101010000000011110010101110010;
		correct = 32'b10111001001110111101000110101111;
		#400 //4.562506e-30 * -3.925874e+25 = -0.00017911823
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010011010111001010111100111010;
		b = 32'b11101101101111100000001010111010;
		correct = 32'b11000001101000111100110001100111;
		#400 //2.7854297e-27 * -7.350681e+27 = -20.474806
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110000001001010100001011001111;
		b = 32'b10101000001000011111000001000010;
		correct = 32'b11011000110100010001010000111011;
		#400 //2.0458317e+29 * -8.989393e-15 = -1839078600000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010001011001101101010100100110;
		b = 32'b00101100111000100000110010111010;
		correct = 32'b10111110110010111101001110100101;
		#400 //-61963657000.0 * 6.4247193e-12 = -0.3980991
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101100111000110110111001111000;
		b = 32'b11110000000100000110100100110011;
		correct = 32'b01011101100000000100101110011001;
		#400 //-6.4639925e-12 * -1.7877208e+29 = 1.1555814e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001011011101110001101111110111;
		b = 32'b01110100001011111110011001010011;
		correct = 32'b01000000001010011100101001110001;
		#400 //4.7591508e-32 * 5.574484e+31 = 2.652981
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010010000001100100000111111011;
		b = 32'b11001111000101111110110101100100;
		correct = 32'b01100001100111110101101011010101;
		#400 //-144158150000.0 * -2548917200.0 = 3.6744718e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100010011001001010011100010000;
		b = 32'b01101100101111001111100010001010;
		correct = 32'b11001111101010001100100010101101;
		#400 //-3.0988204e-18 * 1.827614e+27 = -5663447600.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110010010111110001111011100000;
		b = 32'b10100000011111110110110101111001;
		correct = 32'b10010011010111101001111100101011;
		#400 //1.29873285e-08 * -2.1635562e-19 = -2.8098815e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000001100110011111111010101110;
		b = 32'b10101110001011010010101000001011;
		correct = 32'b00110000010100000101010011001100;
		#400 //-19.249355 * -3.9372988e-11 = 7.5790463e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000011000011000111101000001110;
		b = 32'b11110111001001010011011100110010;
		correct = 32'b01111010101101010101000111101001;
		#400 //-140.47678 * -3.3509706e+33 = 4.7073353e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010000110001011100100010100011;
		b = 32'b11001110100111111001100101111100;
		correct = 32'b11011111111101101001110001100100;
		#400 //26546084000.0 * -1338818000.0 = -3.5540376e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110110101010100001100101010100;
		b = 32'b00110100101111000110000001111010;
		correct = 32'b11101011111110100101010101101000;
		#400 //-1.7250082e+33 * 3.5087925e-07 = -6.0526955e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001000110001110110010010110111;
		b = 32'b01000011000110000101000010001101;
		correct = 32'b10001100011011010100010100010100;
		#400 //-1.2000555e-33 * 152.31465 = -1.8278603e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100000101000100001011011011000;
		b = 32'b01010100100100011110110001110101;
		correct = 32'b01110101101110001100100101001111;
		#400 //9.343808e+19 * 5013899000000.0 = 4.684891e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010001110111001111001101100100;
		b = 32'b11111100111111010001010110111001;
		correct = 32'b01001111010110100110111101001001;
		#400 //-3.485988e-28 * -1.05127335e+37 = 3664726300.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110000110011100000011110011000;
		b = 32'b10011100101110011010000111010110;
		correct = 32'b10001110000101010110010110111100;
		#400 //1.4990631e-09 * -1.2284107e-21 = -1.8414651e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000101000000110001101010100001;
		b = 32'b10000011011011001100001100011100;
		correct = 32'b00001000111100101000000011110000;
		#400 //-2097.6643 * -6.957814e-37 = 1.4595158e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011000010010101000010100011000;
		b = 32'b10101011111011011111101111110001;
		correct = 32'b10000100101111000100010010000110;
		#400 //2.6175083e-24 * -1.6909791e-12 = -4.4261516e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010000111100011001111010001101;
		b = 32'b01001000011111110110011000111101;
		correct = 32'b10011001111100010000110101101101;
		#400 //-9.5302025e-29 * 261528.95 = -2.4924239e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000110000100011011001011111001;
		b = 32'b00111101011100001010111011010010;
		correct = 32'b00000100000010001111101101001001;
		#400 //2.7402957e-35 * 0.05876047 = 1.6102108e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101011000101100011101001010010;
		b = 32'b00010111011010100011110010010010;
		correct = 32'b00000011000010010111010011011010;
		#400 //5.337164e-13 * 7.568593e-25 = 4.039482e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011101100100001010100100000011;
		b = 32'b11000110111000100011101100100001;
		correct = 32'b10100100111111111010110100111100;
		#400 //3.8291237e-21 * -28957.564 = -1.1088209e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000110011111000000110011100001;
		b = 32'b00100010100111000111010000010000;
		correct = 32'b00101001100110100000101000011111;
		#400 //16131.22 * 4.240677e-18 = 6.8407296e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111111001010111000011000101010;
		b = 32'b11110000111010100000101001111010;
		correct = 32'b01110000100111001100111110100111;
		#400 //-0.67001593 * -5.7945726e+29 = 3.882456e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001101110010110000000001011111;
		b = 32'b11110110110100111101100000111100;
		correct = 32'b11000101001001111111110011000110;
		#400 //1.251093e-30 * -2.1483601e+33 = -2687.7983
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000011100111000111001100001111;
		b = 32'b01100101110001011111000000010010;
		correct = 32'b00101001111100011110111010000011;
		#400 //9.195272e-37 * 1.1684184e+23 = 1.0743925e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001110100100011001100011000000;
		b = 32'b11100011010010100101011111110100;
		correct = 32'b01110010011001100010100100011010;
		#400 //-1221353500.0 * -3.73258e+21 = 4.5587994e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100000100100111010110100110001;
		b = 32'b01100100111100110010111110010010;
		correct = 32'b01000110000011000100100011010111;
		#400 //2.5017377e-19 * 3.5887893e+22 = 8978.21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000111101100100011001111100101;
		b = 32'b00100001110110100011000010101011;
		correct = 32'b10101010000101111110001000010010;
		#400 //-91239.79 * 1.4785137e-18 = -1.3489928e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011100011010000001101100000111;
		b = 32'b10001100011100010011011100100011;
		correct = 32'b00101001010110101011001101101111;
		#400 //-2.6132765e+17 * -1.8582557e-31 = 4.8561358e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001001000011110010111100010010;
		b = 32'b11000001101010000111001001010001;
		correct = 32'b01001011001111000110110110101000;
		#400 //-586481.1 * -21.055819 = 12348840.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010101111100100000000001111100;
		b = 32'b01110000001000110010011000010111;
		correct = 32'b01000110100110100011101001010001;
		#400 //9.7743786e-26 * 2.0196842e+29 = 19741.158
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000101100101100011011001011101;
		b = 32'b11001000100110010111100010111110;
		correct = 32'b11001110101101000001101010101101;
		#400 //4806.7954 * -314309.94 = -1510823600.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011110011010110110100011100010;
		b = 32'b00110110111001000010001110101111;
		correct = 32'b00010101110100011100101000111010;
		#400 //1.2462486e-20 * 6.7990836e-06 = 8.4733485e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000111001111101110111111111111;
		b = 32'b00111110110010010000000101000110;
		correct = 32'b11000110100101011110101101100010;
		#400 //-48879.996 * 0.39258784 = -19189.691
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010001010101110100011001100010;
		b = 32'b00011001111000010011010010011111;
		correct = 32'b00101011101111010110000100011100;
		#400 //57787425000.0 * 2.3285708e-23 = 1.3456211e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001000110011010111010010101110;
		b = 32'b10011000000001110110010011101100;
		correct = 32'b10100001010110010101001100001101;
		#400 //420773.44 * -1.7499294e-24 = -7.3632377e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010011001100100010110001111011;
		b = 32'b11000110101010011111111010011011;
		correct = 32'b01011010011011001010000100100010;
		#400 //-765250440000.0 * -21759.303 = 1.6651315e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000001110000011111110111111011;
		b = 32'b11101111100000110011100110010111;
		correct = 32'b10110001110001101110000100110111;
		#400 //7.1261447e-38 * -8.122432e+28 = -5.7881624e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111110001111111001101101010011;
		b = 32'b00010101000110101110000111100101;
		correct = 32'b11010011111001111101100100000110;
		#400 //-6.367226e+37 * 3.1278252e-26 = -1991557000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101001110111100000101010001011;
		b = 32'b10100110100000111110111000000011;
		correct = 32'b10010000111001001101101110101011;
		#400 //9.8606094e-14 * -9.154464e-16 = -9.0268595e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010101111111000111110000011101;
		b = 32'b01101010100000000100110100111000;
		correct = 32'b11000000111111010001010001101110;
		#400 //-1.01977806e-25 * 7.755358e+25 = -7.908744
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110111101010110111010001100000;
		b = 32'b11011001110110010011111011100111;
		correct = 32'b11010010000100010111111111000110;
		#400 //2.043898e-05 * -7643654000000000.0 = -156228490000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111010100111101101011100110000;
		b = 32'b00011110001110101110111001000001;
		correct = 32'b11011001011001111111100001011011;
		#400 //-4.123737e+35 * 9.896028e-21 = -4080861800000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011100110010001100111011000110;
		b = 32'b00110101001111111010001011111010;
		correct = 32'b00010010100101100101001000011101;
		#400 //1.3288339e-21 * 7.1390207e-07 = 9.486573e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100111011011110101101000111000;
		b = 32'b10011100011010010101100011010110;
		correct = 32'b10000100010110100010110000101100;
		#400 //3.321682e-15 * -7.720805e-22 = -2.564606e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000101010111111001001111110111;
		b = 32'b11101011011110100100000100100001;
		correct = 32'b11110001010110101000111101100001;
		#400 //3577.2478 * -3.0253902e+26 = -1.0822571e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011011100101010001011111110111;
		b = 32'b01010101110001110100001100001101;
		correct = 32'b01110001111010000001100101011100;
		#400 //8.393224e+16 * 27386350000000.0 = 2.2985978e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100101010111110011110001101001;
		b = 32'b01011000011101001111011011000110;
		correct = 32'b00111110010101011001110011000101;
		#400 //1.9362635e-16 * 1077362900000000.0 = 0.20860584
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101000101011001010001101100111;
		b = 32'b00000000011010000001110011001110;
		correct = 32'b00101001100011000110101110011101;
		#400 //6.52209e+24 * 9.561225e-39 = 6.235917e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011100111010101100011000000000;
		b = 32'b01000100000100010111100100100011;
		correct = 32'b01100001100001010110100100111110;
		#400 //5.286628e+17 * 581.89276 = 3.0762506e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011111010111010001011001111011;
		b = 32'b10110000000000111011101100110000;
		correct = 32'b00001111111000111000100001010100;
		#400 //-4.6817166e-20 * -4.792353e-10 = 2.243644e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111111011110110010010011101010;
		b = 32'b11111100000110101000000100100010;
		correct = 32'b01111100000101111001001011100100;
		#400 //-0.981032 * -3.2089314e+36 = 3.1480645e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000011111101010110101011011000;
		b = 32'b01010000000010010100011010001001;
		correct = 32'b00010100100000111001100111001100;
		#400 //1.4424336e-36 * 9212405000.0 = 1.3288282e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000000001101010000011010110101;
		b = 32'b11110111100101110110010111100011;
		correct = 32'b11111000010101100001111000000010;
		#400 //2.8285344 * -6.141432e+33 = -1.7371252e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100110000100110011110011000000;
		b = 32'b01001001101000110111010110100000;
		correct = 32'b01110000001111000000011010101010;
		#400 //1.7382713e+23 * 1339060.0 = 2.3276495e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001010011001010000001001100100;
		b = 32'b10111100101100010111001101001011;
		correct = 32'b11000111100111101011110111001010;
		#400 //3752089.0 * -0.021661421 = -81275.58
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110111110001110100011101010000;
		b = 32'b00100000001110010100001110010100;
		correct = 32'b00011000100100000011011100100100;
		#400 //2.3755856e-05 * 1.5692469e-19 = 3.7278805e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011011101111101111000000110110;
		b = 32'b00111001110110101010111100111110;
		correct = 32'b10010110001000110001101101000010;
		#400 //-3.1588096e-22 * 0.00041710766 = -1.3175636e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100100001110100111101011110010;
		b = 32'b11100101111100001101100111011101;
		correct = 32'b11001010101011110111000111110110;
		#400 //4.043646e-17 * -1.4217335e+23 = -5748987.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100100000101011000101001101101;
		b = 32'b10111100100010011001010110000001;
		correct = 32'b10100001001000001011110011010011;
		#400 //3.2426476e-17 * -0.016794922 = -5.4460015e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111111001100001111101110100;
		b = 32'b00110001101010111111011100010111;
		correct = 32'b10101010000110101001010100100000;
		#400 //-2.7432783e-05 * 5.004846e-09 = -1.3729686e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001010001111111000010101111000;
		b = 32'b00110011100100011101000010100100;
		correct = 32'b00111110010110100010110101100000;
		#400 //3137886.0 * 6.79004e-08 = 0.21306372
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011111010101011010000001011010;
		b = 32'b11000010101010110101100101010110;
		correct = 32'b11100010100011101111110010101001;
		#400 //1.5393402e+19 * -85.674484 = -1.3188219e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000100101100001110111011010100;
		b = 32'b01110011010101011100010100100111;
		correct = 32'b10111000100100111011111011111001;
		#400 //-4.159673e-36 * 1.6936614e+31 = -7.045078e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111001110111110100111100110000;
		b = 32'b00001100110011101011110110101001;
		correct = 32'b01000111001101000101011100101010;
		#400 //1.4493604e+35 * 3.1853473e-31 = 46167.164
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010011011010001101001011111110;
		b = 32'b10000101011010100111101010100000;
		correct = 32'b00011001010101010100000001100010;
		#400 //-999972300000.0 * -1.102515e-35 = 1.1024844e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101010000000000000011001101010;
		b = 32'b10110110011101101111010001001110;
		correct = 32'b01100000111101110000000010101110;
		#400 //-3.86932e+25 * -3.679906e-06 = 1.4238734e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101001001110111011100110010010;
		b = 32'b01010010111011111100100010001100;
		correct = 32'b10111100101011111101010101001111;
		#400 //-4.1683298e-14 * 514930900000.0 = -0.021464018
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000010111111100001010011100000;
		b = 32'b10001110100011011111111001101001;
		correct = 32'b10010010000011001110111000000000;
		#400 //127.04077 * -3.500417e-30 = -4.446957e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100100011110111100100010011011;
		b = 32'b00011100110110100011000101111111;
		correct = 32'b00000001110101101001100110000010;
		#400 //5.459687e-17 * 1.4438824e-21 = 7.883146e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111111000011100101000111010100;
		b = 32'b11001001100000011011100101110110;
		correct = 32'b01001001000100000011110010101101;
		#400 //-0.5559361 * -1062702.8 = 590794.8
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100101110010100111110001111101;
		b = 32'b11101010101111100000011110000010;
		correct = 32'b01010001000101100100111001010101;
		#400 //-3.512577e-16 * -1.1486568e+26 = 40347455000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000001001001111011000110010011;
		b = 32'b11001101101000100100010100001000;
		correct = 32'b01001111010101001001011100101110;
		#400 //-10.480853 * -340304130.0 = 3566677500.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101100110100001000101101100111;
		b = 32'b10001101100000010000010110101001;
		correct = 32'b10111010110100100011010110110111;
		#400 //2.016919e+27 * -7.951601e-31 = -0.0016037737
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011010011101011111100000011100;
		b = 32'b01010000000100111101001000100101;
		correct = 32'b01101011000011100000011101100001;
		#400 //1.7308542e+16 * 9920091000.0 = 1.7170231e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000011010011010000101100111001;
		b = 32'b01001001100101110101010011001000;
		correct = 32'b11001101011100100110101100001101;
		#400 //-205.04384 * 1239705.0 = -254193870.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110111111100000001101100111110;
		b = 32'b10010110110010101100101010011011;
		correct = 32'b10001111001111100011001110000110;
		#400 //2.8622915e-05 * -3.2762722e-25 = -9.377646e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101000011010111010110110001001;
		b = 32'b01000101101010111000101001010110;
		correct = 32'b00101110100111011110110001000101;
		#400 //1.308275e-14 * 5489.292 = 7.181503e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111000001000100000000010110011;
		b = 32'b10010101110001101110000101100010;
		correct = 32'b00001110011110111011011001010110;
		#400 //-3.862446e-05 * -8.0327155e-26 = 3.102593e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001000000000010000111011011111;
		b = 32'b10100101111111011001101110110011;
		correct = 32'b00101110011111111011010001100001;
		#400 //-132155.48 * -4.399401e-16 = 5.8140496e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111100010111011100001100111;
		b = 32'b00101101101000011011001001001011;
		correct = 32'b00110101101100001000000010010000;
		#400 //71536.805 * 1.8382759e-11 = 1.3150438e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011011011110110000010100100101;
		b = 32'b00111010100010010001100001101100;
		correct = 32'b00010110100001100110110110110011;
		#400 //2.0763896e-22 * 0.0010459549 = 2.1718098e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001110001110110110111011101010;
		b = 32'b10001011110001100011110011000000;
		correct = 32'b10011010100100010010010001000100;
		#400 //786152060.0 * -7.635823e-32 = -6.0029185e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111111010110101000001001011;
		b = 32'b00001110010010000000100011110101;
		correct = 32'b10000110101101111101111011110110;
		#400 //-2.8051572e-05 * 2.4656216e-30 = -6.916456e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001000110001010000001101001100;
		b = 32'b11100001111110100001111010000100;
		correct = 32'b10101011010000000111110010110100;
		#400 //1.1857281e-33 * -5.767356e+20 = -6.8385163e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100111101100001101110011100011;
		b = 32'b10110001010001100000110100101010;
		correct = 32'b00011001100010001101001111110000;
		#400 //-4.90893e-15 * -2.8820275e-09 = 1.4147671e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111000010111000110010011100111;
		b = 32'b01111101100001010001001001001110;
		correct = 32'b11110110011001010010000001011101;
		#400 //-5.254606e-05 * 2.2110296e+37 = -1.161809e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100010100101010000111100100011;
		b = 32'b10011000000111011011010111100001;
		correct = 32'b10111011001101111010100001011110;
		#400 //1.3748278e+21 * -2.03836e-24 = -0.0028023939
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001011010100100001111100000101;
		b = 32'b11101011111010001101111101000100;
		correct = 32'b10110111101111110010001101011101;
		#400 //4.0467865e-32 * -5.6305026e+26 = -2.2785442e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101010000110010111111111010101;
		b = 32'b11010001111000001010110001101100;
		correct = 32'b00111100100001101011011100111101;
		#400 //-1.363348e-13 * -120620680000.0 = 0.016444797
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010011110100011000101100010001;
		b = 32'b00110111010100111111010001111001;
		correct = 32'b11001011101011010111110110111011;
		#400 //-1799962600000.0 * 1.2633501e-05 = -22739830.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110111001101100100000100010001;
		b = 32'b10001011010001110100000011001000;
		correct = 32'b01000011000011011101101010110011;
		#400 //-3.6965536e+33 * -3.8374742e-32 = 141.8543
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011101010000100011000100000111;
		b = 32'b10010000101100011101111110010001;
		correct = 32'b10101110100001101110110101111101;
		#400 //8.745608e+17 * -7.015865e-29 = -6.135801e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101001010101010010000000010101;
		b = 32'b01111000110111000010100110010101;
		correct = 32'b11100010101101110100101000110000;
		#400 //-4.7323328e-14 * 3.5723397e+34 = -1.69055e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111001001000110000001101010001;
		b = 32'b00011011000110000110011001100011;
		correct = 32'b11010100110000100001011001010101;
		#400 //-5.290073e+34 * 1.2606228e-22 = -6668786600000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010110010010000101000001100101;
		b = 32'b01100001100011101000001111110001;
		correct = 32'b01111000010111110000011110101011;
		#400 //55061904000000.0 * 3.2861813e+20 = 1.809434e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011110101110110010111101100110;
		b = 32'b00110111000000011011110011001111;
		correct = 32'b11010110001111011011100111100001;
		#400 //-6.744056e+18 * 7.73296e-06 = -52151510000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001011110001110111001101001100;
		b = 32'b11110100100000011010010010000000;
		correct = 32'b01000000110010100000001010000110;
		#400 //-7.682549e-32 * -8.217075e+31 = 6.312808
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110010001000111000111001000110;
		b = 32'b11110101111101111110100010011000;
		correct = 32'b01101000100111100110001011100000;
		#400 //-9.520198e-09 * -6.285229e+32 = 5.9836626e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101001000011101010111000101011;
		b = 32'b11000011011000101001010100101111;
		correct = 32'b11101100111111001001000111001111;
		#400 //1.0780622e+25 * -226.58275 = -2.442703e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111100001011101001101000111101;
		b = 32'b01010111010000011111101111010011;
		correct = 32'b11010100000001000100111000001001;
		#400 //-0.01065689 * 213287320000000.0 = -2272979600000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010110111100100001000001011010;
		b = 32'b10111010011110000000001100011110;
		correct = 32'b01010001111010101000001011001010;
		#400 //-133076020000000.0 * -0.0009460914 = 125902080000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101111101011110011010111100011;
		b = 32'b10100111101001100110101110111000;
		correct = 32'b11010111111000111100110101010101;
		#400 //1.0845004e+29 * -4.6191044e-15 = -500942070000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010000111110111100011000111111;
		b = 32'b11001110111101111110110001010010;
		correct = 32'b00100000011100111101010010110010;
		#400 //-9.930749e-29 * -2079729900.0 = 2.0653276e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001101000011000100111011011000;
		b = 32'b10101000110000001001001110011010;
		correct = 32'b00110110010100110001100000001111;
		#400 //-147123580.0 * -2.1380294e-14 = 3.1455454e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000001101011110101110101111011;
		b = 32'b01000101010011001001101010001110;
		correct = 32'b00000111100011000010100001011110;
		#400 //6.4418985e-38 * 3273.6597 = 2.1088584e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011010110111111001011001110;
		b = 32'b00101010001010100110000101110100;
		correct = 32'b10110110000100100110001011110111;
		#400 //-14414542.0 * 1.5132844e-13 = -2.18133e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110001101101100101011011100000;
		b = 32'b11010111000001111001010011101111;
		correct = 32'b11001001010000010010001111001001;
		#400 //5.3067737e-09 * -149073730000000.0 = -791100.56
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110000010000011101011111111011;
		b = 32'b11010100111101010001001110100101;
		correct = 32'b11000101101110011001001010010011;
		#400 //7.051992e-10 * -8420772500000.0 = -5938.322
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001011010011011101111000001111;
		b = 32'b11101000110010010011101000111000;
		correct = 32'b00110100101000011101001000101011;
		#400 //-3.9648622e-32 * -7.602157e+24 = 3.0141504e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011101101001100011111110111110;
		b = 32'b10011110100010010010100010010100;
		correct = 32'b10111100101100100010010011101110;
		#400 //1.4974378e+18 * -1.4522222e-20 = -0.021746125
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110011011000001100001111010010;
		b = 32'b01011110111000101011000110000101;
		correct = 32'b11010010110001110000100010111100;
		#400 //-5.233216e-08 * 8.167492e+18 = -427422500000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111001101111000110110010000101;
		b = 32'b10000110101100010001101010101100;
		correct = 32'b11000001000000100101101010101010;
		#400 //1.2229411e+35 * -6.661919e-35 = -8.147135
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101011011110000100001111101110;
		b = 32'b11000011000101011000000111100111;
		correct = 32'b00101111000100001111110110000100;
		#400 //-8.820157e-13 * -149.50743 = 1.318679e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110001001110100101111110111110;
		b = 32'b10011011001001100011001010101000;
		correct = 32'b01001100111100011111110111101100;
		#400 //-9.228793e+29 * -1.3747566e-22 = 126873440.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000100111001001011111111101101;
		b = 32'b10110101101011010011000000000001;
		correct = 32'b00111011000110101100000010011000;
		#400 //-1829.9977 * -1.2903475e-06 = 0.002361333
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011011100001011010010011100011;
		b = 32'b11101000000100110111000001001000;
		correct = 32'b11000100000110011111000010011000;
		#400 //2.210956e-22 * -2.7850364e+24 = -615.7593
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011100010101110110010100100010;
		b = 32'b10010000001110101101001001011100;
		correct = 32'b10101101000111010011000001111001;
		#400 //2.4251327e+17 * -3.6844087e-29 = -8.93518e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011110010001001111011010111011;
		b = 32'b00101001111011001011010010100100;
		correct = 32'b10001000101101100001111001110000;
		#400 //-1.0427176e-20 * 1.05118415e-13 = -1.0960882e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111101001001011000110010110;
		b = 32'b10110001000011111010001010001010;
		correct = 32'b00101001001110001100111110001000;
		#400 //-1.9633018e-05 * -2.0901632e-09 = 4.1036212e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010011110000101100111011111101;
		b = 32'b10100110110011010011101101110100;
		correct = 32'b00111011000111000010110011111111;
		#400 //-1673392700000.0 * -1.4240847e-15 = 0.002383053
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010100010101100100010100100100;
		b = 32'b00101011100110000010100011000100;
		correct = 32'b11000000011111101011011001011000;
		#400 //-3681132000000.0 * 1.0811564e-12 = -3.9798794
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101111111110100001110101010110;
		b = 32'b11111010011110011000000101101000;
		correct = 32'b11101010111100111100010011110111;
		#400 //4.549558e-10 * -3.2387665e+35 = -1.4734956e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000001000100100101010011100111;
		b = 32'b00110100000111100010111010011011;
		correct = 32'b00110101101101001101011000010101;
		#400 //9.145728 * 1.4731852e-07 = 1.3473351e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010011010110010011100001100010;
		b = 32'b00111101000100111010001101010111;
		correct = 32'b00010000111110101000101111110010;
		#400 //2.741705e-27 * 0.036044445 = 9.8823233e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101010001011000110110100010100;
		b = 32'b10101111000111111110110110011100;
		correct = 32'b10011001110101110110111110010011;
		#400 //1.5314513e-13 * -1.4545382e-10 = -2.2275543e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111100011101101110100100110101;
		b = 32'b00100111100010110111101111100100;
		correct = 32'b11100100100001101000100000011110;
		#400 //-5.12814e+36 * 3.8714573e-15 = -1.9853376e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101011111111100000100001101101;
		b = 32'b00101010101101000011110000000001;
		correct = 32'b00010111001100101101100101111000;
		#400 //1.8050124e-12 * 3.201606e-13 = 5.7789386e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010001100101101001000100101111;
		b = 32'b00001101011010101101100010110011;
		correct = 32'b10011111100010100010000000101001;
		#400 //-80835110000.0 * 7.236766e-31 = -5.849848e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010011100111001110100011110110;
		b = 32'b11101010101011100100000111000000;
		correct = 32'b01111110110101011001110101001000;
		#400 //-1347846700000.0 * -1.0533179e+26 = 1.4197111e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111001101110011100101101100110;
		b = 32'b10110111000011010001010000101000;
		correct = 32'b01110001010011001100011101010000;
		#400 //-1.2058754e+35 * -8.408948e-06 = 1.0140143e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011111011000000001101100100010;
		b = 32'b01110100001111111011100101001000;
		correct = 32'b01010100001001111101011001110001;
		#400 //4.745629e-20 * 6.0759683e+31 = 2883429000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100000111100011110010111100101;
		b = 32'b11011001010011100111100100010100;
		correct = 32'b11111010110000110001100101100111;
		#400 //1.3944472e+20 * -3632310800000000.0 = -5.0650655e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110111001111100001001100100000;
		b = 32'b00101110010100001111010000011000;
		correct = 32'b01100110000110110010010011000110;
		#400 //3.855173e+33 * 4.7510523e-11 = 1.8316129e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011101010101101000010010000000;
		b = 32'b10100001000110010100011100001000;
		correct = 32'b00111111000000000111000010110110;
		#400 //-9.661013e+17 * -5.1932425e-19 = 0.50171983
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011111000110010011011000111011;
		b = 32'b00101011001000101110110001001111;
		correct = 32'b10001010110000110000001101111101;
		#400 //-3.244387e-20 * 5.7881906e-13 = -1.8779129e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111101010110010100101010001011;
		b = 32'b00111000110011001100110100000000;
		correct = 32'b10110110101011011101010101100111;
		#400 //-0.053049605 * 9.765662e-05 = -5.180645e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111111101001000011011111101100;
		b = 32'b10011001100000010001101110110100;
		correct = 32'b10011001101001011010001111100111;
		#400 //1.2829566 * -1.3349477e-23 = -1.71268e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011100000101111000000100000011;
		b = 32'b10111010111101010001000110010101;
		correct = 32'b11010111100100010000100011100000;
		#400 //1.7057829e+17 * -0.0018697256 = -318934600000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001011000110001111011001000110;
		b = 32'b00000101010001000110011100110111;
		correct = 32'b00010000111010101011010001110011;
		#400 //10024518.0 * 9.234833e-36 = 9.257475e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001100001110010100111000101110;
		b = 32'b11011010010010011111011010001001;
		correct = 32'b10100111000100100011000011010110;
		#400 //1.4275408e-31 * -1.4211885e+16 = -2.0288044e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011100111010011011111100010010;
		b = 32'b10111111000101010010101011111001;
		correct = 32'b00011100100010000011001101110010;
		#400 //-1.5468037e-21 * -0.58268696 = 9.013023e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010000100011010000100100101101;
		b = 32'b10000110011011100011111010100111;
		correct = 32'b10010111100000110100000100001100;
		#400 //18929510000.0 * -4.4808855e-35 = -8.482097e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011011000101100100100110100000;
		b = 32'b10110010000111011110001011011001;
		correct = 32'b00001101101110010110000010100111;
		#400 //-1.2431499e-22 * -9.190182e-09 = 1.14247735e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110100000000010110011001101011;
		b = 32'b10100100111010110000000001011110;
		correct = 32'b10011001011011011001001001100111;
		#400 //1.205132e-07 * -1.01915626e-16 = -1.22821785e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100001111100111100101100001010;
		b = 32'b01101110000110000110000001100100;
		correct = 32'b01010000100100010001110001011001;
		#400 //1.6520064e-18 * 1.1789563e+28 = 19476433000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001011001101011010100000110101;
		b = 32'b11010110111001011101001100001001;
		correct = 32'b10100010101000110001010100110111;
		#400 //3.4985877e-32 * -126347280000000.0 = -4.42037e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000001010110100011010101000111;
		b = 32'b10001111100100101000110010011111;
		correct = 32'b10010001011110011101010001111110;
		#400 //13.638007 * -1.4450877e-29 = -1.9708116e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011000001000010001110100101011;
		b = 32'b10010001001001001100000110111011;
		correct = 32'b10101001110011110110000100111000;
		#400 //708586600000000.0 * -1.2997017e-28 = -9.2095114e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110101100011001111110011100111;
		b = 32'b01001010000000110011111101001111;
		correct = 32'b01000000000100001001000010010000;
		#400 //1.0504417e-06 * 2150355.8 = 2.2588234
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110100100100000010000000000011;
		b = 32'b10000110100010010101111001101111;
		correct = 32'b10111011100110101010110010011000;
		#400 //9.13501e+31 * -5.167243e-35 = -0.004720282
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101101110001010111000111100100;
		b = 32'b01011010110100111110011110000010;
		correct = 32'b11001001001000110110111101101101;
		#400 //-2.2446885e-11 * 2.9822883e+16 = -669430.8
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111100101110101010101100100001;
		b = 32'b00101001110110110010110111010101;
		correct = 32'b11100111000111111101000111010001;
		#400 //-7.753905e+36 * 9.733504e-14 = -7.547267e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011001001111011000000011101100;
		b = 32'b10011101010000111101110011101001;
		correct = 32'b10110111000100001111110010111011;
		#400 //3333782600000000.0 * -2.5922243e-21 = -8.641912e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100001101100010101001101111011;
		b = 32'b00110000110111101101111010000010;
		correct = 32'b00010011000110100110000010000101;
		#400 //1.2016084e-18 * 1.6215866e-09 = 1.948512e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011110111110010011010000011011;
		b = 32'b01001101111011111111010000011011;
		correct = 32'b11101101011010011001010101000101;
		#400 //-8.9785037e+18 * 503219040.0 = -4.518154e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111000001001000000101011111;
		b = 32'b00110100111001001000001111111010;
		correct = 32'b00111100011011001000111100010000;
		#400 //33921.37 * 4.2564335e-07 = 0.014438406
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001110011010111110110011001111;
		b = 32'b00001100010001111100100110001001;
		correct = 32'b10011011001110000001111011010000;
		#400 //-989541300.0 * 1.539105e-31 = -1.5230079e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101000010111100001000101001011;
		b = 32'b11010100011010100010010101100000;
		correct = 32'b00111101010010110001110000111010;
		#400 //-1.2327225e-14 * -4022597600000.0 = 0.049587466
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111101011010001100010010010111;
		b = 32'b11001011001100100110010111010111;
		correct = 32'b01001001001000100011010101001010;
		#400 //-0.056828108 * -11691479.0 = 664404.6
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001000111000001001100100000100;
		b = 32'b11011111011000000101010110110100;
		correct = 32'b00101000110001001101000100010100;
		#400 //-1.3517483e-33 * -1.6165024e+19 = 2.1851044e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001100110110010111100110101111;
		b = 32'b00000110000001110110110011111111;
		correct = 32'b10010011011001100001011110000110;
		#400 //-114019704.0 * 2.5470756e-35 = -2.904168e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011111111111100101011100110000;
		b = 32'b00111011011011011111000010010011;
		correct = 32'b00011011111011000110010110111011;
		#400 //1.07717424e-19 * 0.0036306723 = 3.9108667e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111010010010001001010010000;
		b = 32'b11011011011100001110011100000000;
		correct = 32'b11100011001111010011011011010111;
		#400 //51474.562 * -6.780798e+16 = -3.4903863e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000110001101001010011101100101;
		b = 32'b00110011111110100100011011111110;
		correct = 32'b10111010101100001001110110010010;
		#400 //-11561.849 * 1.16544456e-07 = -0.0013474694
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000101110100010010101000111101;
		b = 32'b11001011010101100001001111101101;
		correct = 32'b10010001101011101110100110010111;
		#400 //1.9669781e-35 * -14029805.0 = -2.759632e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010111011001000010011110000;
		b = 32'b11000110111110001010000111110001;
		correct = 32'b01000010011001011011011001100111;
		#400 //-0.001804499 * -31824.97 = 57.428127
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100010001010001011100000100001;
		b = 32'b01111010010111101110011001111111;
		correct = 32'b11011101000100101110011110010110;
		#400 //-2.2865723e-18 * 2.8934123e+35 = -6.6159965e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010101100010010101101001110010;
		b = 32'b11000111101110010111000101110111;
		correct = 32'b01011101110001101111111001111010;
		#400 //-18877694000000.0 * -94946.93 = 1.792379e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100010110000110000010101000111;
		b = 32'b10011001110001011001110000011101;
		correct = 32'b10111101000101101000100111111101;
		#400 //1.7987477e+21 * -2.0432376e-23 = -0.03675269
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101101111110001111000011111000;
		b = 32'b10101100000011111100100011001001;
		correct = 32'b10011010100010111101000111011010;
		#400 //2.8301347e-11 * -2.043298e-12 = -5.7828086e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001010100011110010000111001100;
		b = 32'b00011001000100010000000100010111;
		correct = 32'b10100100001000100010010110000001;
		#400 //-4690150.0 * 7.496544e-24 = -3.5159917e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111001101010001101101111010000;
		b = 32'b00010101010101101001011010001111;
		correct = 32'b01001111100011011000101100001111;
		#400 //1.0959552e+35 * 4.3335726e-26 = 4749401600.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111011101101100001001000001;
		b = 32'b01110011011011101010110101000000;
		correct = 32'b01111011011001100000111110010111;
		#400 //63170.254 * 1.8909921e+31 = 1.1945445e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011100011110100000001111010100;
		b = 32'b11010111110011000111010010011100;
		correct = 32'b01110100110001111010110011101111;
		#400 //-2.8149181e+17 * -449602400000000.0 = 1.265594e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110111101100000011010110111;
		b = 32'b00110100011101010010110011001101;
		correct = 32'b10101011111010111001111101111011;
		#400 //-7.332153e-06 * 2.2833702e-07 = -1.6742019e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111000101011110010101110011011;
		b = 32'b01110111100111000100000100000101;
		correct = 32'b11110000110101011101011000100000;
		#400 //-8.3527724e-05 * 6.3384146e+33 = -5.2943335e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001010011010110101101001000010;
		b = 32'b11111010011111000011100101100011;
		correct = 32'b11000101011001111110000110011011;
		#400 //1.1331814e-32 * -3.2740569e+35 = -3710.1003
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011101010011101001101011110001;
		b = 32'b10000000011111010011110110110110;
		correct = 32'b00011110010010100010011011101011;
		#400 //-9.304673e+17 * -1.1501575e-38 = 1.0701839e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010010000111100100110001110;
		b = 32'b01001011011001101011001100000101;
		correct = 32'b11000110001100000110111111111111;
		#400 //-0.00074686937 * 15119109.0 = -11291.999
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001001010011110011110001000011;
		b = 32'b11001000111100010101101000111000;
		correct = 32'b10010010110000110110000011000100;
		#400 //2.4945054e-33 * -494289.75 = -1.2330085e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111011110101101010110001100110;
		b = 32'b01010110100001001111101000001110;
		correct = 32'b01010010110111110000010100101001;
		#400 //0.006551313 * 73104756000000.0 = 478932140000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110011101010110011010101110000;
		b = 32'b00010000001011001010010011000111;
		correct = 32'b00000100011001101110110000110101;
		#400 //7.972528e-08 * 3.404796e-29 = 2.7144831e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000010000000111110001111000111;
		b = 32'b10111011110100000010001101010101;
		correct = 32'b10111110010101100111011010001011;
		#400 //32.97244 * -0.006351868 = -0.20943658
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101011110100100110110010111101;
		b = 32'b01110010101010000000010001110100;
		correct = 32'b11011111000010100001101100000101;
		#400 //-1.4951578e-12 * 6.655855e+30 = -9.951553e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001010000010101000110010001110;
		b = 32'b11011000100110011011011110001101;
		correct = 32'b11100011001001100110001010101111;
		#400 //2269987.5 * -1352109000000000.0 = -3.0692704e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001011000101100100010001001101;
		b = 32'b10010011010100110000100010001100;
		correct = 32'b10011110111101111011111010100000;
		#400 //9847885.0 * -2.6636158e-27 = -2.6230983e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110011100000010010001001100101;
		b = 32'b10100101001010001000000011010011;
		correct = 32'b01011001001010011111111100011100;
		#400 //-2.0462155e+31 * -1.4615325e-16 = 2990610400000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010000110100000011110000110100;
		b = 32'b00000000000111001001101111010101;
		correct = 32'b10010000101110100010101010111011;
		#400 //-27948851000.0 * 2.627296e-39 = -7.34299e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001010011010110011000011110100;
		b = 32'b10110100111011101111101111101100;
		correct = 32'b00111111110110111000111011110101;
		#400 //-3853373.0 * -4.4514252e-07 = 1.7153002
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011101001101110000000000001111;
		b = 32'b11000111111000101101000100110010;
		correct = 32'b10100101101000100010001110011000;
		#400 //2.4219879e-21 * -116130.39 = -2.812664e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000000001100101000010110000;
		b = 32'b11000100101100111101011110010010;
		correct = 32'b00110101001111001011011100001011;
		#400 //-4.886358e-10 * -1438.7366 = 7.030182e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110110000001000111011000101010;
		b = 32'b00110101011000001111011101000111;
		correct = 32'b11101011111010001100111010101111;
		#400 //-6.7166e+32 * 8.380634e-07 = -5.6289365e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001000000110000111011101000100;
		b = 32'b10010011000100100111101011110100;
		correct = 32'b10011011101011100111101001111110;
		#400 //156125.06 * -1.8488411e-27 = -2.8865044e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001000111111011001101111000111;
		b = 32'b11000110001000101101011001001000;
		correct = 32'b10001111101000010101000011011011;
		#400 //1.5263507e-33 * -10421.57 = -1.590697e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111100000111100010011000110101;
		b = 32'b01011111010110010101001101101100;
		correct = 32'b11011100000001100100000111101100;
		#400 //-0.009652664 * 1.5659979e+19 = -1.5116051e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001001111010000010001011100101;
		b = 32'b11010011100111010111011001111101;
		correct = 32'b11011110000011101100100011011000;
		#400 //1901660.6 * -1352595500000.0 = -2.5721777e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011100001000011110100101001011;
		b = 32'b01011010100101100011011110001010;
		correct = 32'b11110111001111100000001110100101;
		#400 //-1.8229592e+17 * 2.1141156e+16 = -3.8539466e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010010111101100001111111000011;
		b = 32'b11110110101000000111110101001100;
		correct = 32'b01001010000110100100110001010000;
		#400 //-1.55326125e-27 * -1.6275563e+33 = 2528020.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110001010001111110111001001100;
		b = 32'b01000010101110101001111010001011;
		correct = 32'b00110100100100011011111011110101;
		#400 //2.9093767e-09 * 93.309654 = 2.7147294e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011001110010010010011111011000;
		b = 32'b01011111101100011010000111000001;
		correct = 32'b00111010000010111001001110100110;
		#400 //2.0799006e-23 * 2.5599448e+19 = 0.00053244305
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000101101101001110011001001000;
		b = 32'b10010101111010100000101001101001;
		correct = 32'b00011100001001010110000111011001;
		#400 //-5788.785 * -9.452827e-26 = 5.4720386e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111100000111100110010111000000;
		b = 32'b00110110011101101100010000011110;
		correct = 32'b11110011000110001010111100011111;
		#400 //-3.2897866e+36 * 3.6771012e-06 = -1.2096878e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010110010011001101111110100001;
		b = 32'b00111010000001000110111101111100;
		correct = 32'b10010000110100111111100100001110;
		#400 //-1.6549554e-25 * 0.0005052013 = -8.3608555e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010100110001010000111001000001;
		b = 32'b10010100001001001000011101011010;
		correct = 32'b10101001011111010100101010100011;
		#400 //6770781600000.0 * -8.3065775e-27 = -5.6242022e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001001010100111011111111010100;
		b = 32'b10111000111110110111111000011101;
		correct = 32'b10000010110100000000010101100101;
		#400 //2.5488398e-33 * -0.00011992103 = -3.056595e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100110011100100010111010110000;
		b = 32'b01010110110111111000101110010000;
		correct = 32'b11111101110100110111101010110011;
		#400 //-2.8591848e+23 * 122895255000000.0 = -3.5138025e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110001111010100101001001000100;
		b = 32'b10110001010010011010110110010010;
		correct = 32'b00100011101110001001100101110111;
		#400 //-6.819649e-09 * -2.9348013e-09 = 2.0014315e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000000101110010010111011101;
		b = 32'b10111100000011001101100100011010;
		correct = 32'b00101100101001100101000111000111;
		#400 //-5.4987287e-10 * -0.008596683 = 4.727083e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000000101100111010001000000100;
		b = 32'b00111001111111100101000101110011;
		correct = 32'b10111011001100100111001111100111;
		#400 //-5.6135273 * 0.0004850734 = -0.0027229728
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011000011000011111110100011100;
		b = 32'b10101111000000110111111101011111;
		correct = 32'b00000111111010000010100111101100;
		#400 //-2.9208356e-24 * -1.1959632e-10 = 3.493212e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000111101001000000001001001010;
		b = 32'b01101111010010000000010101000001;
		correct = 32'b00110111100000000010010100101000;
		#400 //2.4677323e-34 * 6.1903354e+28 = 1.5276091e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010110110001101101101010011110;
		b = 32'b11110010001010000111101101011110;
		correct = 32'b11001001100000101101111101001100;
		#400 //3.2126592e-25 * -3.337128e+30 = -1072105.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000110100101011101111001001100;
		b = 32'b01011101001111101000111011001110;
		correct = 32'b11100100010111110001110100101101;
		#400 //-19183.148 * 8.581962e+17 = -1.6462905e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001100111110101001100000011010;
		b = 32'b01001011011110011111110101110101;
		correct = 32'b01011000111101001011011000001100;
		#400 //131383500.0 * 16383349.0 = 2152501800000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111110000001100100101111010001;
		b = 32'b01010011111001010001111101000110;
		correct = 32'b11010010011100000110010001110100;
		#400 //-0.13114859 * 1968144400000.0 = -258119370000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000011101100010110000101000010;
		b = 32'b11010011111010011000001111100110;
		correct = 32'b10011000001000011100110011101001;
		#400 //1.0425454e-36 * -2005880500000.0 = -2.0912215e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011001111110111010111011110000;
		b = 32'b10001000001110010110111101001001;
		correct = 32'b00100010101101100100111011010100;
		#400 //-8855320600000000.0 * -5.5802228e-34 = 4.941466e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000111111010101001111000000110;
		b = 32'b11110111101100010010000110111001;
		correct = 32'b11000000001000100101011000101010;
		#400 //3.5301285e-34 * -7.1853166e+33 = -2.536509
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111001010000101100111011111111;
		b = 32'b00001001011110000111111110111010;
		correct = 32'b01000011001111010001100110111001;
		#400 //6.3219e+34 * 2.991197e-33 = 189.10048
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100110101111111111111001101001;
		b = 32'b00011001010001010100110001000010;
		correct = 32'b11000000100100111111011111111000;
		#400 //-4.5333252e+23 * 1.02000614e-23 = -4.6240196
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010110101001101101111011110011;
		b = 32'b01001101100100010100011001000000;
		correct = 32'b00100100101111010110010000100101;
		#400 //2.6959447e-25 * 304662530.0 = 8.2135336e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100110100100111110010001011011;
		b = 32'b01000100001111111011001000110111;
		correct = 32'b11101011010111010111110010101001;
		#400 //-3.4920014e+23 * 766.7846 = -2.677613e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011011011110100001001010101110;
		b = 32'b11011011100011111110010101000100;
		correct = 32'b01110111100011001001000001100100;
		#400 //-7.0389283e+16 * -8.1006e+16 = 5.701954e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001101101010110101110101100111;
		b = 32'b11101100010000010111010011010010;
		correct = 32'b01111010100000010111111110011110;
		#400 //-359378140.0 * -9.354974e+26 = 3.3619734e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100000111111111001110010001001;
		b = 32'b10001110111100001000000101110111;
		correct = 32'b10110000011100000010010000000101;
		#400 //1.4734998e+20 * -5.9289238e-30 = -8.736268e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000101000001111111001101001111;
		b = 32'b10111110000111100001001010111011;
		correct = 32'b01000011101001111110010000111010;
		#400 //-2175.2068 * -0.15436833 = 335.78302
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010101110000110010110001010011;
		b = 32'b00110010110010010001000101111010;
		correct = 32'b11001001000110010100101100100000;
		#400 //-26824392000000.0 * 2.3407427e-08 = -627890.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100101110001101001101001100001;
		b = 32'b00010110100000100101000010101000;
		correct = 32'b10111100110010100011000111110000;
		#400 //-1.1723454e+23 * 2.1053534e-25 = -0.024682015
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011101101000011111110011011101;
		b = 32'b01110011111001110011000111011110;
		correct = 32'b11010010000100100100101010111001;
		#400 //-4.28778e-21 * 3.6634277e+31 = -157079720000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010011001010100110010111111100;
		b = 32'b00101111101100011100011101101111;
		correct = 32'b00000011011011001010101010000101;
		#400 //2.1507299e-27 * 3.2337819e-10 = 6.9549914e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100101001110110001101100110100;
		b = 32'b00111101010110001100001010101010;
		correct = 32'b01100011000111100110110100111011;
		#400 //5.522402e+22 * 0.05292002 = 2.9224564e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001010110111001000000011011010;
		b = 32'b01101001000001000110110001111011;
		correct = 32'b01110100011001000001111111000001;
		#400 //7225453.0 * 1.0005656e+25 = 7.2295394e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011011011101110101100100011001;
		b = 32'b01000010100110100001111001110001;
		correct = 32'b11011110100101001110100100000011;
		#400 //-6.9622283e+16 * 77.059456 = -5.3650554e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111110101011011001010110110110;
		b = 32'b10001000011100110001000111011110;
		correct = 32'b00000111101001001101000100111001;
		#400 //-0.33903283 * -7.3146155e-34 = 2.4798947e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010010101111101000101110011011;
		b = 32'b01010010011011010011100101001111;
		correct = 32'b01100101101100001001000111100110;
		#400 //409193000000.0 * 254717180000.0 = 1.0422848e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111110101010010111000001110010;
		b = 32'b01100111100100001011111110101010;
		correct = 32'b11100110101111111001110000110111;
		#400 //-0.330936 * 1.3671127e+24 = -4.5242683e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101000000010100110000001010001;
		b = 32'b00110111001000111011011000111010;
		correct = 32'b01011111101100001111101110100111;
		#400 //2.6138532e+24 * 9.757985e-06 = 2.550594e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111111011001111001100001001110;
		b = 32'b00110010110101100110011001000110;
		correct = 32'b01110010110000011111010111010111;
		#400 //3.0784248e+38 * 2.4959387e-08 = 7.6835596e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010101110100110100101101010101;
		b = 32'b11011100010111110001101111011101;
		correct = 32'b01110010101110000010010110011110;
		#400 //-29040063000000.0 * -2.5119822e+17 = 7.294812e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100101111101100111111010011101;
		b = 32'b01000001111111010010010111101110;
		correct = 32'b00101000011100111011111110100111;
		#400 //4.2759994e-16 * 31.64352 = 1.3530768e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111101001111010101111001100101;
		b = 32'b00110100000100000011101111101001;
		correct = 32'b00110001110101010110001011010100;
		#400 //0.0462326 * 1.343284e-07 = 6.2103513e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010111001010101011110101100010;
		b = 32'b11011101011000000000101111110011;
		correct = 32'b11110101000101010110110110101110;
		#400 //187730370000000.0 * -1.0090165e+18 = -1.8942305e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011111101001111110001001000011;
		b = 32'b01100001111011001001000101100011;
		correct = 32'b01000010000110110010001111101110;
		#400 //7.110157e-20 * 5.4548848e+20 = 38.785088
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011000101110000000010101111000;
		b = 32'b11011001111111010110101101101110;
		correct = 32'b10110011001101100010101010100001;
		#400 //4.7568407e-24 * -8916411000000000.0 = -4.2413948e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000001100101001111100111000001;
		b = 32'b00111000010000000010111011100100;
		correct = 32'b10111010010111111010110100110101;
		#400 //-18.62195 * 4.5820037e-05 = -0.0008532585
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101010101000100000001101110001;
		b = 32'b01110110000100110010010001110010;
		correct = 32'b01100001001110100011111000010101;
		#400 //2.877937e-13 * 7.461004e+32 = 2.14723e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111100110000001111100101100001;
		b = 32'b00001000110011101111101100100000;
		correct = 32'b11000110000111000000010111111001;
		#400 //-8.015832e+36 * 1.2457213e-33 = -9985.493
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100111101111101010110101100101;
		b = 32'b11010010100001100010011011111100;
		correct = 32'b10111010110001111101011110011001;
		#400 //5.292359e-15 * -288089830000.0 = -0.0015246748
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110000101111110100011101000000;
		b = 32'b10100111100001001100110111001100;
		correct = 32'b10011000110001100111010100000011;
		#400 //1.391733e-09 * -3.6860485e-15 = -5.1299952e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010011001010010101011010111010;
		b = 32'b01000011110101000010010011100000;
		correct = 32'b01010111100011000101010000110110;
		#400 //727304500000.0 * 424.2881 = 308586620000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010111000100001000001011000010;
		b = 32'b00111111110110011110010111001111;
		correct = 32'b01010111011101100000000100100001;
		#400 //158891270000000.0 * 1.7023257 = 270484710000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011011110011001011011010010011;
		b = 32'b01011110101011001001001100101000;
		correct = 32'b01111011000010100000000001011000;
		#400 //1.15243275e+17 * 6.2176635e+18 = 7.165439e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110100011101001000111000011001;
		b = 32'b01000000001111111100001001010101;
		correct = 32'b00110101001101110010111110101010;
		#400 //2.2775966e-07 * 2.996236 = 6.824217e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001010000010001011010010000110;
		b = 32'b11001010111000101011011001011000;
		correct = 32'b10010101011100100010000101111011;
		#400 //6.5821145e-33 * -7428908.0 = -4.8897922e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011100111110110000110000000001;
		b = 32'b11011111011100110110110100100010;
		correct = 32'b11111100111011101011011101101010;
		#400 //5.6530734e+17 * -1.7540714e+19 = -9.915894e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111000101111110001111001010000;
		b = 32'b00110010100000101011101101100000;
		correct = 32'b00101011110000110011001010001111;
		#400 //9.113236e-05 * 1.52192e-08 = 1.3869616e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111001110011111111001010011000;
		b = 32'b10101111100100111101010110111100;
		correct = 32'b00101001111100000010101111010110;
		#400 //-0.00039662863 * -2.6891012e-10 = 1.06657454e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100100000111111001111101001100;
		b = 32'b01001100110001001010001000110110;
		correct = 32'b11110001011101010011011000110101;
		#400 //-1.1778043e+22 * 103092660.0 = -1.21422975e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001011101001110111011011101100;
		b = 32'b01010000110110011011001100011010;
		correct = 32'b01011101000011100110100011110111;
		#400 //21949912.0 * 29219148000.0 = 6.413577e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100111110100111010110111011;
		b = 32'b10111101111100111101010011000101;
		correct = 32'b11000011011011101000110111101011;
		#400 //2003.6791 * -0.11905817 = -238.55437
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011011111100001011001101101011;
		b = 32'b01100100110100010100100000110011;
		correct = 32'b11000001010001001100011001011101;
		#400 //-3.9820616e-22 * 3.0884576e+22 = -12.298429
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111111010010011110010100110000;
		b = 32'b11111001100000101011010000000111;
		correct = 32'b01111001010011100010100010111010;
		#400 //-0.7886534 * -8.483125e+34 = 6.690245e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101011000110001101010101001110;
		b = 32'b10011000000110010111000001001111;
		correct = 32'b11000011101101110011010100010000;
		#400 //1.8476403e+26 * -1.9831488e-24 = -366.41455
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100010001111110010000001110001;
		b = 32'b00110100000110111110111010110001;
		correct = 32'b00010110111010001101010110110001;
		#400 //2.5902501e-18 * 1.4522335e-07 = 3.761648e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100010111110011111001110000011;
		b = 32'b00100111110110001011100101000110;
		correct = 32'b00001011010100111001101001011100;
		#400 //6.7749413e-18 * 6.0152917e-15 = 4.075325e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001101011100101101011001100001;
		b = 32'b00111010101001010111111001111110;
		correct = 32'b01001000100111001111110000101010;
		#400 //254633490.0 * 0.0012626199 = 321505.3
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111011101010000001011111111001;
		b = 32'b00010111111101110101001010011100;
		correct = 32'b00010100001000100110010101011111;
		#400 //0.005129811 * 1.5982854e-24 = 8.198902e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100000000011110011001011011001;
		b = 32'b10100000111001001111110110010101;
		correct = 32'b10000001100000000001011100100010;
		#400 //1.2129395e-19 * -3.879251e-19 = -4.705297e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001101110001000111100111111110;
		b = 32'b01110010011010000000100001011000;
		correct = 32'b01000000101100100001010011110110;
		#400 //1.2108801e-30 * 4.595879e+30 = 5.5650587
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111100010010001001111110001110;
		b = 32'b00100011100011111001111110010100;
		correct = 32'b01100000011000010001110001011111;
		#400 //4.166782e+36 * 1.5571675e-17 = 6.4883778e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100100100110001000000101110110;
		b = 32'b10110101011011110111011110000110;
		correct = 32'b01011010100011101010100000010001;
		#400 //-2.250587e+22 * -8.920837e-07 = 2.0077119e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010010100111100001110001011101;
		b = 32'b01000110111000100011011000101101;
		correct = 32'b00011010000010111011011010000000;
		#400 //9.978194e-28 * 28955.088 = 2.889195e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101011101010101011110010010011;
		b = 32'b00010101011000001111110100010100;
		correct = 32'b11000001100101100000110111001010;
		#400 //-4.128158e+26 * 4.5436083e-26 = -18.756733
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011110110011001100110010001001;
		b = 32'b11001111110100110110101111101010;
		correct = 32'b01101111001010010010001011101010;
		#400 //-7.3786604e+18 * -7094129700.0 = 5.2345175e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100011100000100001011001010;
		b = 32'b10101001110110110000100110001101;
		correct = 32'b10101110110011011001001000011001;
		#400 //961.0436 * -9.7272105e-14 = -9.348273e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010100101100010000011110100100;
		b = 32'b01000000011000110011011001010110;
		correct = 32'b00010101100111010001111101011010;
		#400 //1.7875446e-26 * 3.5501914 = 6.346126e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101111000000000100100110001110;
		b = 32'b10111101101011000011011001011001;
		correct = 32'b00101101001011001001100101001111;
		#400 //-1.1667664e-10 * -0.084088035 = 9.811109e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000011110101001011011001101;
		b = 32'b11001001000000101011010011111111;
		correct = 32'b00111001111111111110001101111111;
		#400 //-9.116377e-10 * -535375.94 = 0.00048806888
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101010001010000101101001001000;
		b = 32'b10101001100001001101100100011011;
		correct = 32'b01010100001011101011101010100111;
		#400 //-5.088147e+25 * -5.8996394e-14 = 3001823300000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111100000100001110100000011110;
		b = 32'b10100011010101101000001011000010;
		correct = 32'b00011111111100101101100000011010;
		#400 //-0.008844404 * -1.1628652e-17 = 1.02848497e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101111111001111010111000110101;
		b = 32'b10011110110000000110011010001010;
		correct = 32'b11001111001011100001111101110100;
		#400 //1.4340328e+29 * -2.03712e-20 = -2921297000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010011100110100100000101111001;
		b = 32'b11101111110000100100101101011000;
		correct = 32'b11000011111010100010011000001000;
		#400 //3.8939626e-27 * -1.2026235e+29 = -468.29712
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000011011010001001011100100101;
		b = 32'b10101010110000111010001111011010;
		correct = 32'b10101110101100011011111111111111;
		#400 //232.59041 * -3.4752653e-13 = -8.0831335e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010101000010001100000010000110;
		b = 32'b00100111100100100100010000110111;
		correct = 32'b10111101000111000100010001111010;
		#400 //-9397529000000.0 * 4.05971e-15 = -0.03815124
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100010101010000111010001100001;
		b = 32'b00011000011100001111100101101011;
		correct = 32'b10111011100111101001000100111011;
		#400 //-1.5537195e+21 * 3.1145197e-24 = -0.00483909
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101000010010010001100110000001;
		b = 32'b00010001101011110111100011010010;
		correct = 32'b10111010100010011101011101011000;
		#400 //-3.7986645e+24 * 2.7684593e-28 = -0.0010516448
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011111010000000010000000011001;
		b = 32'b11101100110111001101011111110110;
		correct = 32'b01001100101001011011110110101001;
		#400 //-4.0684132e-20 * -2.1358682e+27 = 86895944.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011101001001010010010111001101;
		b = 32'b00101011111100011101011100011100;
		correct = 32'b10001001100111000000001101011011;
		#400 //-2.185711e-21 * 1.7183785e-12 = -3.755879e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110001000010111011010010001;
		b = 32'b00000110101101111100110000011010;
		correct = 32'b00000101011001111101100011111001;
		#400 //0.15767886 * 6.913685e-35 = 1.09014194e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110010001010000001011110000000;
		b = 32'b11110111110110110011011000010010;
		correct = 32'b01101010100011111110111110011011;
		#400 //-9.78423e-09 * -8.892263e+33 = 8.700395e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100101000011111011101001101;
		b = 32'b10111100111111111111110011010101;
		correct = 32'b11000010001000011111010101001100;
		#400 //1295.7281 * -0.03124849 = -40.489548
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011011000101010001011111001101;
		b = 32'b00111010101110101011100111111000;
		correct = 32'b11010110010110010111111100110011;
		#400 //-4.196594e+16 * 0.0014246097 = -59785085000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010011001101110000100001111111;
		b = 32'b10001100010001011010010111001101;
		correct = 32'b00100000000011010101000000010101;
		#400 //-786121560000.0 * -1.5226222e-31 = 1.1969661e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001110101011111000010011000110;
		b = 32'b00100101100101110100000011001010;
		correct = 32'b00110100110011110110011101111001;
		#400 //1472357100.0 * 2.6238227e-16 = 3.863204e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001001100001001000110000100000;
		b = 32'b01001000001111110110000101111001;
		correct = 32'b01010010010001100010111000000111;
		#400 //1085828.0 * 195973.89 = 212793930000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100000111110101110010100101001;
		b = 32'b01101001000001100001011011111110;
		correct = 32'b01001010100000110110101001111100;
		#400 //4.2503293e-19 * 1.013154e+25 = 4306238.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111001001101111000110110000111;
		b = 32'b10010000110100010010100001111011;
		correct = 32'b01001010100101011111011110010010;
		#400 //-5.9566303e+34 * -8.2498335e-29 = 4914121.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001000100010001111100010000001;
		b = 32'b00111001000010110001110000100010;
		correct = 32'b11000010000101001101101111110111;
		#400 //-280516.03 * 0.00013266553 = -37.21481
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011110010100101111000010111110;
		b = 32'b10110110000000010000001101000101;
		correct = 32'b01010100110101001001110000000011;
		#400 //-3.7999644e+18 * -1.92244e-06 = 7305204000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111010011101101100111110110010;
		b = 32'b01010001001010001110011101001111;
		correct = 32'b01001100001000101101011101001110;
		#400 //0.0009415104 * 45339700000.0 = 42687800.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000101010010100001011100011011;
		b = 32'b01101000000011110100000101001111;
		correct = 32'b10101101111000100010110011101101;
		#400 //-9.502238e-36 * 2.7060126e+24 = -2.5713176e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111111011110010100111001110101;
		b = 32'b10000101011100100000101001000010;
		correct = 32'b10000101011010111011011000101000;
		#400 //0.9738534 * -1.13806694e-35 = -1.1083104e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010100000111111110011101000110;
		b = 32'b00111000100111011100101110101011;
		correct = 32'b10001101010001010010000000011010;
		#400 //-8.073059e-27 * 7.5242795e-05 = -6.0743953e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101010000010100000111011101010;
		b = 32'b10110111011100101011100010110101;
		correct = 32'b00100010000000101110010110110110;
		#400 //-1.2262037e-13 * -1.44673295e-05 = 1.7739893e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100001011001100100101100110101;
		b = 32'b01011100111100000010011110011011;
		correct = 32'b01111110110110000000101000100011;
		#400 //2.6551065e+20 * 5.4078033e+17 = 1.4358294e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111011101011011010110111100;
		b = 32'b01011100001100001110000101010110;
		correct = 32'b11010100001010011100010100111001;
		#400 //-1.4645451e-05 * 1.9914942e+17 = -2916633300000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001110010010100111111100010011;
		b = 32'b01101011000001001111011001110100;
		correct = 32'b10111001110100100101100011101111;
		#400 //-2.4959606e-30 * 1.6074205e+26 = -0.00040120582
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100011100101011100001110100100;
		b = 32'b01111100101000001011011000011100;
		correct = 32'b01100000101111000000100110100000;
		#400 //1.623747e-17 * 6.675689e+36 = 1.08396295e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011111110000101000111110101100;
		b = 32'b11011010001110100000100000110101;
		correct = 32'b10111010100011010110001010100000;
		#400 //8.239988e-20 * -1.3090842e+16 = -0.0010786839
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110010100011010000010010110111;
		b = 32'b00000000001001111110010110011011;
		correct = 32'b10110010101011111101000110010100;
		#400 //-5.586315e+30 * 3.663951e-39 = -2.0467986e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111100101110011010111011010101;
		b = 32'b11101011000110111000010000100001;
		correct = 32'b01101000011000011001100101100010;
		#400 //-0.022666374 * -1.8800746e+26 = 4.2614475e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101001111101101010010001100101;
		b = 32'b00100001100011001101110111110010;
		correct = 32'b01001100000001111011011110111100;
		#400 //3.727151e+25 * 9.545517e-19 = 35577584.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010010101101000110111110111100;
		b = 32'b11100001111000101101001111110001;
		correct = 32'b00110101000111111110000000000110;
		#400 //-1.1387142e-27 * -5.2302952e+20 = 5.955811e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010101100101011010001001010100;
		b = 32'b01001101010000100010111010110100;
		correct = 32'b10100011011000110000000010100000;
		#400 //-6.043673e-26 * 203615040.0 = -1.2305827e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010110110110001100001100000001;
		b = 32'b00010010010001100111011110000100;
		correct = 32'b10101001101010000000110000000101;
		#400 //-119166020000000.0 * 6.26251e-28 = -7.462784e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000101101111011010100101000100;
		b = 32'b00001100111100001001111101111010;
		correct = 32'b10010011001100100100010011010110;
		#400 //-6069.158 * 3.7073836e-31 = -2.2500697e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011011001110011111001010100;
		b = 32'b10000000001001001110110010000010;
		correct = 32'b00001011100001010110100110011011;
		#400 //-15154772.0 * -3.390921e-39 = 5.1388634e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111011111000111010000010100100;
		b = 32'b10111001101001100000000101100110;
		correct = 32'b01110110000100111001101101101001;
		#400 //-2.3638191e+36 * -0.0003166303 = 7.484568e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111001001100001011010011001010;
		b = 32'b00100010011000111011101011110001;
		correct = 32'b00011100000111010011000101011001;
		#400 //0.00016852017 * 3.0863203e-18 = 5.2010723e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110110110010111000111011010;
		b = 32'b11100010110101101010011000101000;
		correct = 32'b01011010001101100101001001001110;
		#400 //-6.480358e-06 * -1.979788e+21 = 1.2829735e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100110111000001101101110011010;
		b = 32'b10110100111101010100000010010001;
		correct = 32'b10011100010101110110101011100001;
		#400 //1.5602645e-15 * -4.5681784e-07 = -7.127567e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010110100011011010000101001101;
		b = 32'b01000110110111101011001110010001;
		correct = 32'b10011101111101100110101001110010;
		#400 //-2.2881574e-25 * 28505.783 = -6.522572e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010000100100011001110110010111;
		b = 32'b00111010001001001011101011010100;
		correct = 32'b01001011001110110110011001110100;
		#400 //19544193000.0 * 0.0006283943 = 12281460.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010100101101100110011001100011;
		b = 32'b00100000010000111010101011000111;
		correct = 32'b00110101100010110110100110101011;
		#400 //6267214500000.0 * 1.6573648e-19 = 1.038706e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011100000011011111000110011101;
		b = 32'b10011101011000011001110010001001;
		correct = 32'b00111001111110100011000001001100;
		#400 //-1.5981451e+17 * -2.9859429e-21 = 0.000477197
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011100011001001101110111011111;
		b = 32'b01000001100100010111111001000100;
		correct = 32'b00011110100000100001001010001101;
		#400 //7.5725634e-22 * 18.186653 = 1.3771958e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010011110100010011011100000000;
		b = 32'b11001010011100001101110000010110;
		correct = 32'b11011110110001001101011101101101;
		#400 //1797141800000.0 * -3946245.5 = -7.0919627e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011100001100111111011100011110;
		b = 32'b00111111111011011000101010100110;
		correct = 32'b11011100101001101111110100111111;
		#400 //-2.0262292e+17 * 1.8557937 = -3.7602635e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001011010001010011000001011001;
		b = 32'b01001101011101110101110001001011;
		correct = 32'b01011001001111101000100010111101;
		#400 //12922969.0 * 259376300.0 = 3351912000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111101001101001010001111110111;
		b = 32'b11100101011000001111001011100001;
		correct = 32'b11100011000111101011101011011010;
		#400 //0.04410168 * -6.639315e+22 = -2.9280496e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010101110011110011011101101000;
		b = 32'b11001001100010000001000000001111;
		correct = 32'b00011111110111000100010011011110;
		#400 //-8.369405e-26 * -1114625.9 = 9.3287555e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110100000101000001101011000011;
		b = 32'b11101100110001110000011110101100;
		correct = 32'b01100001011001100100101001111100;
		#400 //-1.379331e-07 * -1.9248997e+27 = 2.655074e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001001011110111100001001011111;
		b = 32'b11010000111101010110010111101011;
		correct = 32'b10011010111100010101010101000000;
		#400 //3.0304419e-33 * -32936778000.0 = -9.981299e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100101100101011101010000000001;
		b = 32'b01000011111011111100110011111110;
		correct = 32'b01101010000011000101100011100111;
		#400 //8.844292e+22 * 479.6015 = 4.241736e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100101011001011010001010111001;
		b = 32'b10101101000111111110011011010011;
		correct = 32'b01010011000011110110111100011110;
		#400 //-6.7776477e+22 * -9.089357e-12 = 616044560000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001110100000111111100101110110;
		b = 32'b10101101001001000110011010110000;
		correct = 32'b00111100001010011000000101111111;
		#400 //-1107082000.0 * -9.345122e-12 = 0.010345816
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000110001001001001110101001011;
		b = 32'b00101101111010111110100100101110;
		correct = 32'b00110100100101111011001001010101;
		#400 //10535.323 * 2.681996e-11 = 2.8255695e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011100011000101111011111001010;
		b = 32'b01000111100010001100110010010101;
		correct = 32'b10100100011100101001001000001010;
		#400 //-7.5097387e-22 * 70041.164 = -5.2599085e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000010011100110011011111110101;
		b = 32'b00011010001110010101111111111100;
		correct = 32'b00011101001100000001111010100001;
		#400 //60.804646 * 3.833464e-23 = 2.330924e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101001101100111001000010110011;
		b = 32'b11111010011010101111111110100101;
		correct = 32'b11100100101001001101010110010100;
		#400 //7.974298e-14 * -3.0504564e+35 = -2.4325248e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101100001000100001101011111111;
		b = 32'b01000001111110101100001101011110;
		correct = 32'b01101110100111101100101000010011;
		#400 //7.838939e+26 * 31.345394 = 2.4571462e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111110001111101000010110011010;
		b = 32'b00010011001100101100110100110010;
		correct = 32'b01010010000001010001000110011011;
		#400 //6.3311755e+37 * 2.2567928e-27 = 142881500000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010100110010011000011001111101;
		b = 32'b11010011011110000011110111010001;
		correct = 32'b11101000110000110110101011110011;
		#400 //6924358000000.0 * -1066189000000.0 = -7.3826746e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001010000000011011000101000110;
		b = 32'b11001011101101101000011111001010;
		correct = 32'b10010110001110001111000110100101;
		#400 //6.2444655e-33 * -23924628.0 = -1.4939651e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111000111000000001110101001000;
		b = 32'b01001011011000100110100001100101;
		correct = 32'b01000100110001100011010100111110;
		#400 //0.000106866064 * 14837861.0 = 1585.6638
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111100010101111111111000010000;
		b = 32'b00000000011100101110110110000011;
		correct = 32'b00111101010000011110111100010000;
		#400 //4.4859873e+36 * 1.055445e-38 = 0.04734713
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100110100001111110010101000100;
		b = 32'b00010111001110111100100111110110;
		correct = 32'b00111110010001110101111101011101;
		#400 //3.2087434e+23 * 6.067787e-25 = 0.19469972
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101100100011111100101001100111;
		b = 32'b10011101100100001011011010100010;
		correct = 32'b10001010101000101001000011011110;
		#400 //4.0867756e-12 * -3.830532e-21 = -1.5654526e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101010001000011100100100010001;
		b = 32'b10110111011001100010111111001110;
		correct = 32'b11100010000100010111100011011011;
		#400 //4.889664e+25 * -1.3720199e-05 = -6.708716e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010100000101010101001110011;
		b = 32'b01011000111001100000111000010100;
		correct = 32'b11010011111010101101100010100110;
		#400 //-0.0009969011 * 2023585100000000.0 = -2017314200000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111110011011000110011000111010;
		b = 32'b00000101110101011111100101100111;
		correct = 32'b11000100110001011001011101011101;
		#400 //-7.855715e+37 * 2.012204e-35 = -1580.7301
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001110110110010011110101010100;
		b = 32'b10110000011010000101111100110010;
		correct = 32'b00111111110001010011000001011100;
		#400 //-1822337500.0 * -8.453639e-10 = 1.5405383
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011000111010100010101010001000;
		b = 32'b11110011100000011001110000001101;
		correct = 32'b11001100111011010001110001011001;
		#400 //6.0530528e-24 * -2.0537457e+31 = -124314310.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001001000100101100111100000000;
		b = 32'b11111011001000100101000100101001;
		correct = 32'b11000100101110100010101100010010;
		#400 //1.7671442e-33 * -8.427982e+35 = -1489.346
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010001001110100000001111111001;
		b = 32'b00100111010110000100110100000101;
		correct = 32'b10111001000111010010101101010001;
		#400 //-49933160000.0 * 3.0017774e-15 = -0.00014988823
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010101110011000011011010000111;
		b = 32'b00000001011101001111011110001001;
		correct = 32'b00010111110000110110100101101111;
		#400 //28066820000000.0 * 4.499332e-38 = 1.2628195e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010111110110100110100100010111;
		b = 32'b01111011101001010000111101011000;
		correct = 32'b01010100000011001101001011010011;
		#400 //1.4114448e-24 * 1.7140804e+36 = 2419329900000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000000001111100000101101010000;
		b = 32'b10111100001101110111100101001010;
		correct = 32'b10111101000010000011010000100000;
		#400 //2.9694405 * -0.011198351 = -0.033252835
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101001100110101100000100110011;
		b = 32'b11111011100110001000110111111110;
		correct = 32'b11100101101110000111000100011000;
		#400 //6.8724886e-14 * -1.5842181e+36 = -1.0887521e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011011110001011011010010110;
		b = 32'b10011010011010011100101100010001;
		correct = 32'b00100110011000110010001101111000;
		#400 //-16299670.0 * -4.8347306e-23 = 7.8804515e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011010000101011111011010000001;
		b = 32'b10101110111100010001100000101100;
		correct = 32'b11001001100011010011101100111000;
		#400 //1.0552701e+16 * -1.0963705e-10 = -1156967.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011010001101100100010010000001;
		b = 32'b11000111011101000000000001111111;
		correct = 32'b01100010001011011011100110100101;
		#400 //-1.2825942e+16 * -62464.496 = 8.0116596e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100001110111110011100110011110;
		b = 32'b10110000001111001110101100110101;
		correct = 32'b10010010101001001011101101101000;
		#400 //1.5126319e-18 * -6.872825e-10 = -1.0396054e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010001100010010011011011011101;
		b = 32'b11011001001000111100000110101001;
		correct = 32'b11101011001011111000101101110111;
		#400 //73666370000.0 * -2880834500000000.0 = -2.1222062e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011111101101010100111110001010;
		b = 32'b10011110000111100111101011111010;
		correct = 32'b00111110011000000111110001100000;
		#400 //-2.6129626e+19 * -8.389881e-21 = 0.21922445
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110100100010111111011000000100;
		b = 32'b10010111101010010100110000110001;
		correct = 32'b00001100101110010001111000100001;
		#400 //-2.6069768e-07 * -1.0940602e-24 = 2.8521896e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010111001110100011110000000010;
		b = 32'b11110011111000010111000000100110;
		correct = 32'b11001011101001000000000001010100;
		#400 //6.017558e-25 * -3.572209e+31 = -21495976.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101011101011011111000010000000;
		b = 32'b00100011011010111001101001110111;
		correct = 32'b10001111101000000001010010111001;
		#400 //-1.2359141e-12 * 1.2772085e-17 = -1.57852e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110010001000100000100001100;
		b = 32'b10000100100010111001001001001001;
		correct = 32'b10000011010101011111111011101101;
		#400 //0.19165438 * -3.2813085e-36 = -6.2887715e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000110100001101110101100100101;
		b = 32'b01000111100100011111001100001101;
		correct = 32'b11001110100110011101011010010000;
		#400 //-17269.572 * 74726.1 = -1290487800.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101011100110110011001001101100;
		b = 32'b00110111000111111100101010000110;
		correct = 32'b00100011010000011011111000110000;
		#400 //1.1027407e-12 * 9.524292e-06 = 1.0502825e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100111111100101100110000101001;
		b = 32'b11000101000111001000100011011111;
		correct = 32'b10101101100101000111011000111001;
		#400 //6.7389844e-15 * -2504.5544 = -1.6878153e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000111010111001100111011111111;
		b = 32'b00000110001110010000111111011011;
		correct = 32'b10001110000111111001111101000011;
		#400 //-56526.996 * 3.4806282e-35 = -1.9674945e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110011010011111010011101010110;
		b = 32'b01100010000101011000000110100111;
		correct = 32'b11010101111100101000101100100000;
		#400 //-4.8348134e-08 * 6.894768e+20 = -33334919000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111110001010101110010111000110;
		b = 32'b00000001111010110100110001111010;
		correct = 32'b11000000100111010001001111111010;
		#400 //-5.6790453e+37 * 8.6435105e-38 = -4.9086885
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000010000110100100101010001110;
		b = 32'b11011111101111000010011110001011;
		correct = 32'b00100010011000101100110100101011;
		#400 //-1.1335529e-37 * -2.7115916e+19 = 3.0737326e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011110111110111001000111101011;
		b = 32'b10110110100001100111011110010010;
		correct = 32'b00010110000001000010001111100001;
		#400 //-2.6636009e-20 * -4.007431e-06 = 1.0674196e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100001101000101110001110011101;
		b = 32'b00010001110100100101111000100001;
		correct = 32'b00110100000001011101101010011011;
		#400 //3.7559673e+20 * 3.319017e-28 = 1.2466118e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110011101100001001000000000100;
		b = 32'b10010111011010001101001010000011;
		correct = 32'b00001011101000001001001110110100;
		#400 //-8.221835e-08 * -7.5228946e-25 = 6.1852e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011111101101100101100111001100;
		b = 32'b00010110010001010011111110011101;
		correct = 32'b00110110100011001000000001101010;
		#400 //2.6279515e+19 * 1.5933606e-25 = 4.1872745e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010000001101000101000101101001;
		b = 32'b10000010001101111101110110110101;
		correct = 32'b10010011000000011000001001011100;
		#400 //12100937000.0 * -1.3508343e-37 = -1.6346361e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101010001101110001000100100100;
		b = 32'b10100100110000100010111011100110;
		correct = 32'b01001111100010101101110010000111;
		#400 //-5.5328592e+25 * -8.421354e-17 = 4659416600.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011110111101011100100001101111;
		b = 32'b01011000110000011011100001101000;
		correct = 32'b01111000001110011111110100101000;
		#400 //8.855264e+18 * 1703982100000000.0 = 1.5089212e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100110011001110111001000101101;
		b = 32'b00111010001010110111101101010001;
		correct = 32'b01100001000110110000100011000001;
		#400 //2.732432e+23 * 0.0006541508 = 1.7874226e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010111001111011101000101001100;
		b = 32'b00110100010110001101000010011110;
		correct = 32'b11001100001000001100001101000111;
		#400 //-208706620000000.0 * 2.0192462e-07 = -42143004.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010110011010011111110011110000;
		b = 32'b10101111111111011000001100101000;
		correct = 32'b10000110111001111011011011011010;
		#400 //1.8901403e-25 * -4.6113624e-10 = -8.716122e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110011000011001101100010000101;
		b = 32'b11001000001001101000011010000000;
		correct = 32'b00111011101101110011110011001100;
		#400 //-3.2793213e-08 * -170522.0 = 0.0055919643
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011011101010101100100000011011;
		b = 32'b01001011110111111010100110110011;
		correct = 32'b10101000000101010011010110000101;
		#400 //-2.8253456e-22 * 29315942.0 = -8.282767e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011010100000110111101111111001;
		b = 32'b00101000010100001011101010111110;
		correct = 32'b10000011010101100110100101001000;
		#400 //-5.438062e-23 * 1.1586813e-14 = -6.3009805e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011000000001111000000100000110;
		b = 32'b00110110011101010010100110100010;
		correct = 32'b00001111000000011100010010000100;
		#400 //1.7513481e-24 * 3.6532078e-06 = 6.3980386e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001111100111001101011101110010;
		b = 32'b01001110001010111100100010010101;
		correct = 32'b00011110010100100111110110011010;
		#400 //1.5465774e-29 * 720512300.0 = 1.1143281e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100001111100010011101000010011;
		b = 32'b00001000100111111111011010101100;
		correct = 32'b10101011000101101011101110000010;
		#400 //-5.5623125e+20 * 9.627457e-34 = -5.3550925e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111110001110101000100011100010;
		b = 32'b00110011011111011000001000000011;
		correct = 32'b10110010001110001011100000000011;
		#400 //-0.18216279 * 5.9024398e-08 = -1.0752049e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101010001000010011100111010111;
		b = 32'b01011101011010010101001000101110;
		correct = 32'b11001000000100101111000101100110;
		#400 //-1.431974e-13 * 1.0507844e+18 = -150469.6
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000110000111101101111001011;
		b = 32'b00100111110001011110110100011011;
		correct = 32'b10011001000101110110110110001010;
		#400 //-1.4250586e-09 * 5.4935554e-15 = -7.828638e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001101111000101010011101100001;
		b = 32'b00000011010011110010010100011100;
		correct = 32'b10010001101101110110011000110010;
		#400 //-475327520.0 * 6.087443e-37 = -2.8935292e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111101111111111011010000010100;
		b = 32'b01110001111110010010010100000011;
		correct = 32'b11110000011110001101101100011111;
		#400 //-0.12485519 * 2.4674084e+30 = -3.0806873e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111101001000111111011000001110;
		b = 32'b10011011111100111101011101000111;
		correct = 32'b11011001100111000010110001110000;
		#400 //1.362136e+37 * -4.0340097e-22 = -5494869500000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011001100000001010001110000100;
		b = 32'b00111110000110110110000000110001;
		correct = 32'b11011000000111000010011010101110;
		#400 //-4526073000000000.0 * 0.15173413 = -686759800000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011111011101001111011101000110;
		b = 32'b10001001111111111100100101101010;
		correct = 32'b00101001111101001100001100001010;
		#400 //-1.7651654e+19 * -6.1578426e-33 = 1.08696106e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011101111101110101111000101000;
		b = 32'b11111111010000010010010110001001;
		correct = 32'b11011101101110101010001001000001;
		#400 //6.547771e-21 * -2.567359e+38 = -1.6810479e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001110110010101001111110000011;
		b = 32'b11101110110110000101011111001011;
		correct = 32'b10111110001010110011110000010011;
		#400 //4.995045e-30 * -3.3477449e+28 = -0.16722135
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110011111010000110000100101110;
		b = 32'b01000000001010000010111000011100;
		correct = 32'b11110100100110001010100110100001;
		#400 //-3.6822019e+31 * 2.6278143 = -9.676143e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100111100101000100110010111011;
		b = 32'b11001111011100000001110100101100;
		correct = 32'b10110111100010110001100011010101;
		#400 //4.1161443e-15 * -4028443600.0 = -1.6581655e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110010100010000111011000000;
		b = 32'b11011111100111000100110101001010;
		correct = 32'b01010110011111110100100000110110;
		#400 //-3.1152013e-06 * -2.252548e+19 = 70171402000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001000100011101111010000101001;
		b = 32'b01100001100110001011010011101011;
		correct = 32'b00101010101010101000101111111110;
		#400 //8.603716e-34 * 3.521177e+20 = 3.0295205e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011110110011101100010100010101;
		b = 32'b01111110110101011001000001110110;
		correct = 32'b11011110001011000111111010101001;
		#400 //-2.189261e-20 * 1.4193782e+38 = -3.1073895e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111000100101111001010011101101;
		b = 32'b10101000101001000100001001101111;
		correct = 32'b11100001110000101000010101111100;
		#400 //2.4595544e+34 * -1.8236469e-14 = -4.4853586e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001110100010011100011101010011;
		b = 32'b10110110110111010100001101100110;
		correct = 32'b00000101111011100010101010110001;
		#400 //-3.396505e-30 * -6.5941595e-06 = 2.2397095e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011101011100111000011100101000;
		b = 32'b01100000110110010011001100111100;
		correct = 32'b01111110110011101001111001001110;
		#400 //1.0967524e+18 * 1.2520735e+20 = 1.3732147e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011100111110010110010011110111;
		b = 32'b11000111000001100111000000001111;
		correct = 32'b00100100100000101111100000000100;
		#400 //-1.6503537e-21 * -34416.06 = 5.679867e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001100000010110111110110111001;
		b = 32'b00111101011111111001110110000100;
		correct = 32'b00001010000010110100100000001111;
		#400 //1.0746004e-31 * 0.062406078 = 6.706159e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001110010010100010000101011010;
		b = 32'b01101110010110000010001111011010;
		correct = 32'b00111101001010101010100001110011;
		#400 //2.491448e-30 * 1.6723026e+28 = 0.041664552
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110100011011011101100011100010;
		b = 32'b10010111110100000110100010111001;
		correct = 32'b01001100110000011010000110000100;
		#400 //-7.5376786e+31 * -1.3468121e-24 = 101518370.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000000110110110100110000111;
		b = 32'b10010011001101110011000000010110;
		correct = 32'b00000011110111100110101101000001;
		#400 //-5.6538635e-10 * -2.3121556e-27 = 1.3072612e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110010000010111100001101010111;
		b = 32'b11111000011110100110001001000000;
		correct = 32'b11101011000010001011001001100111;
		#400 //8.13528e-09 * -2.0313546e+34 = -1.652564e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100000111001111010101011000101;
		b = 32'b11011010000000011010101110101100;
		correct = 32'b10111011011010101011000011010000;
		#400 //3.9245928e-19 * -9124757000000000.0 = -0.0035810955
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111100101101010110100110111000;
		b = 32'b10110011100011011011110100111010;
		correct = 32'b11110000110010001110001010100101;
		#400 //7.5356e+36 * -6.600244e-08 = -4.97368e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001100010110111011001011001100;
		b = 32'b11000000000000001101011010100110;
		correct = 32'b01001100110111010010001100111000;
		#400 //-57592624.0 * -2.013101 = 115939780.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010100111100011100110110001010;
		b = 32'b10001011100011101111111111010101;
		correct = 32'b10100001000001110001000110100111;
		#400 //8308284000000.0 * -5.5081344e-32 = -4.576314e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000010110010110010010011101101;
		b = 32'b00110110001011100010011010011000;
		correct = 32'b00111001100010100011000110111001;
		#400 //101.57212 * 2.5950485e-06 = 0.00026358457
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111011001110001010101001000111;
		b = 32'b01011100001111010010010100110101;
		correct = 32'b11011000000010000111000010001101;
		#400 //-0.0028177665 * 2.1295872e+17 = -600067900000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100111111110011001010001101011;
		b = 32'b00001000100011111101000000010100;
		correct = 32'b10110001000011000011010011000100;
		#400 //-2.3572142e+24 * 8.655418e-34 = -2.0402675e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110011011111100001011100100101;
		b = 32'b01000101010010101101000111111111;
		correct = 32'b10111001010010010100111010110001;
		#400 //-5.9160033e-08 * 3245.1248 = -0.00019198169
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001001100000110110000101001001;
		b = 32'b11001001100110101111111011110111;
		correct = 32'b10010011100111110001011010111110;
		#400 //3.162859e-33 * -1269726.9 = -4.015967e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110010011011111100101000111000;
		b = 32'b11000010111000111001000110000010;
		correct = 32'b11110101110101010010100010011011;
		#400 //4.7495286e+30 * -113.784195 = -5.404213e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011100101000001001101000001;
		b = 32'b10100101100111010111011111100010;
		correct = 32'b00110001101101100010101001001101;
		#400 //-19408514.0 * -2.7316394e-16 = 5.301706e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000000011100101011001001010010;
		b = 32'b01000011000100110001010001110100;
		correct = 32'b10000100000000111100101100011110;
		#400 //-1.0533216e-38 * 147.0799 = -1.5492243e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001011010011011110100111110100;
		b = 32'b01011010010000101100101111101001;
		correct = 32'b00100110000111001010111101001111;
		#400 //3.965757e-32 * 1.3707587e+16 = 5.436096e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001001011101000001000001110001;
		b = 32'b11000101111000110010011110100111;
		correct = 32'b11001111110110001001000001100010;
		#400 //999687.06 * -7268.9565 = -7266682000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010000001011000010001111001101;
		b = 32'b10011111101100011011111011110110;
		correct = 32'b10110000011011110000101001010001;
		#400 //11552110000.0 * -7.5278334e-20 = -8.6962354e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010000011010001101110110110100;
		b = 32'b00111101110110101100000001111000;
		correct = 32'b11001110110001101111101111011111;
		#400 //-15627375000.0 * 0.10681242 = -1669197700.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001101010000001111001110000100;
		b = 32'b11101101011110011001100101011110;
		correct = 32'b10111011001111000010000001110100;
		#400 //5.945769e-31 * -4.8279486e+27 = -0.0028705867
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101111000111111000001101001010;
		b = 32'b11001100101111110010100011101000;
		correct = 32'b00111100011011100011100011100011;
		#400 //-1.4507609e-10 * -100222780.0 = 0.01453993
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101110000000010100010011001001;
		b = 32'b10100110001000001001100000000111;
		correct = 32'b11010100101000100010111110000100;
		#400 //1.0001681e+28 * -5.5717187e-16 = -5572655000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001110000111000111001100110011;
		b = 32'b11100000110001011000001101011100;
		correct = 32'b11101111011100010110100111011011;
		#400 //656198850.0 * -1.1385856e+20 = -7.471386e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110000100010101000111101010101;
		b = 32'b10011001001100001101100110010111;
		correct = 32'b11001010001111110111000010011111;
		#400 //3.4305767e+29 * -9.142929e-24 = -3136551.8
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001001100101101110110101100100;
		b = 32'b01110010100001111101101111111010;
		correct = 32'b11111100101000000011000111000000;
		#400 //-1236396.5 * 5.3819407e+30 = -6.6542124e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011001111011011100100010101101;
		b = 32'b10110000001101011100111011101101;
		correct = 32'b10001010101010001101111100010110;
		#400 //2.4586278e-23 * -6.6141476e-10 = -1.6261727e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111100000110001011011001010100;
		b = 32'b00101011001001100111010010000101;
		correct = 32'b10100111110001101001011101111001;
		#400 //-0.009320814 * 5.913675e-13 = -5.5120267e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010011010001110010010110011101;
		b = 32'b11101011001101011000110100010000;
		correct = 32'b11111111000011010011101101010100;
		#400 //855329540000.0 * -2.1948172e+26 = -1.877292e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010001110010111101010001000111;
		b = 32'b10100010010100011001100001101010;
		correct = 32'b10110100101001101110000110101000;
		#400 //109429970000.0 * -2.840547e-18 = -3.1084096e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011111100010001010001010010101;
		b = 32'b10111111010110010101011010010101;
		correct = 32'b01011111011010000000000000001101;
		#400 //-1.9691191e+19 * -0.8489774 = 1.6717376e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100010011001001100001100010110;
		b = 32'b00011110111000011000011010001100;
		correct = 32'b11000001110010011000011110110010;
		#400 //-1.0549788e+21 * 2.3878449e-20 = -25.191257
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011100011100101011101111100001;
		b = 32'b10000011001100000011101011111101;
		correct = 32'b00100000001001110001100100011001;
		#400 //-2.7329408e+17 * -5.1789467e-37 = 1.4153754e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100110011111000001100100011101;
		b = 32'b10001101110011010111110110010001;
		correct = 32'b00110100110010100101101111000011;
		#400 //-2.976249e+23 * -1.2664329e-30 = 3.7692197e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011111101001111000100100101001;
		b = 32'b00100001011101100011010011001100;
		correct = 32'b00000001101000010010000001011011;
		#400 //7.0954164e-20 * 8.341792e-19 = 5.918849e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100101011001101100101111101000;
		b = 32'b11000100110101011011110000100111;
		correct = 32'b11101010110000001011000101001001;
		#400 //6.8119106e+22 * -1709.8798 = -1.1647548e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111010111010011100000011011111;
		b = 32'b10111101010011100101101011111001;
		correct = 32'b11111000101111000110110001000101;
		#400 //6.0685853e+35 * -0.050379727 = -3.0573368e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010000011000101000000011100101;
		b = 32'b00100011100101110011111011101010;
		correct = 32'b10110100100001011101000110110001;
		#400 //-15200392000.0 * 1.6398098e-17 = -2.492575e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110101101110100110110001010001;
		b = 32'b10011011110000010101010111010011;
		correct = 32'b11010010000011001100101000101001;
		#400 //4.7263874e+32 * -3.1984634e-22 = -151171780000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110010111101000100001010010100;
		b = 32'b00111011111000101001101100010100;
		correct = 32'b00101111010110000011011010111110;
		#400 //2.8435615e-08 * 0.0069154594 = 1.9664534e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110101000000111000101011101101;
		b = 32'b10010011110011011000101000111111;
		correct = 32'b00001001010100110011101010010010;
		#400 //-4.9003467e-07 * -5.1885597e-27 = 2.542574e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010101000100110100010100011110;
		b = 32'b01010101100000000011000000110010;
		correct = 32'b10101011000100110111110010010001;
		#400 //-2.9740937e-26 * 17618060000000.0 = -5.239776e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011110110011001100010000010101;
		b = 32'b10101001011110101000010111000001;
		correct = 32'b01001000110010000110001001111001;
		#400 //-7.3774707e+18 * -5.5627164e-14 = 410387.78
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111100010111000101100100001101;
		b = 32'b00011010111000100100111011110010;
		correct = 32'b11010111110000101100101010010001;
		#400 //-4.576446e+36 * 9.359895e-23 = -428350540000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001111110100111100001011010010;
		b = 32'b01101001101100111101000100100010;
		correct = 32'b11111010000101001011111000110111;
		#400 //-7105520600.0 * 2.7173165e+25 = -1.9307949e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011010100100110111111101011111;
		b = 32'b00010100111010110110010111010101;
		correct = 32'b00110000000001111010000010011000;
		#400 //2.0758434e+16 * 2.3769102e-26 = 4.934093e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011111010100000011000110001000;
		b = 32'b00001010111000010010001111101101;
		correct = 32'b00101010101101110001100011000000;
		#400 //1.5001921e+19 * 2.1680226e-32 = 3.2524504e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001001010101000010101110111011;
		b = 32'b00111010000010011001100000100011;
		correct = 32'b01000011111001000001001011111100;
		#400 //869051.7 * 0.00052488054 = 456.14832
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011010011011100000100010110101;
		b = 32'b00101111011000110011111011001010;
		correct = 32'b00001010010100110100110000011010;
		#400 //4.922428e-23 * 2.0667837e-10 = 1.01735936e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101000111010011100000010011111;
		b = 32'b01001001101100000010101001101110;
		correct = 32'b00110011001000001101101100101011;
		#400 //2.5951733e-14 * 1443149.8 = 3.7452235e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100110111101111101100110001001;
		b = 32'b01001110100101000011010000111001;
		correct = 32'b01110110000011110111110001010011;
		#400 //5.8521867e+23 * 1243225200.0 = 7.275586e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111110000000000110100010111001;
		b = 32'b10110010111001111000100010111110;
		correct = 32'b00110001011010000100011000101100;
		#400 //-0.12539949 * -2.6954122e-08 = 3.3800331e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111110011101111101011011000;
		b = 32'b01100111000100110011101101000010;
		correct = 32'b01101111011011100001001111100110;
		#400 //105973.69 * 6.95281e+23 = 7.368149e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011101010111001111110100100111;
		b = 32'b01010000110011111110100110011100;
		correct = 32'b01101110101100110111101001011100;
		#400 //9.952454e+17 * 27905548000.0 = 2.777287e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100100011010010011110011101010;
		b = 32'b00111101010000111011001011100011;
		correct = 32'b10100010001100100100110001100001;
		#400 //-5.0575417e-17 * 0.04777802 = -2.4163933e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111011000100101111110111000010;
		b = 32'b00111100000000000101100100100110;
		correct = 32'b11110111100100110110010000100010;
		#400 //-7.632222e+35 * 0.007833755 = -5.978895e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010110000111111100011010100101;
		b = 32'b01110000110010010111101100100000;
		correct = 32'b11000111011110110111111110100000;
		#400 //-1.2906599e-25 * 4.988427e+29 = -64383.625
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111001010101000010100001011100;
		b = 32'b00110010000111110111101110011011;
		correct = 32'b00101100000001000010101110000001;
		#400 //0.0002023293 * 9.283123e-09 = 1.8782478e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111100111110001110010000110100;
		b = 32'b11010000110011101011010100000110;
		correct = 32'b11001110010010001111011110100001;
		#400 //0.030382253 * -27743760000.0 = -842917950.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111010101100110110011000011001;
		b = 32'b00101111010110100010100101011111;
		correct = 32'b11101010100110001110000111101111;
		#400 //-4.6574596e+35 * 1.9841682e-10 = -9.241183e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111111100010110100000001000101;
		b = 32'b10101000010000101100111000101111;
		correct = 32'b00101000010100111110110110110111;
		#400 //-1.0878989 * -1.0813872e-14 = 1.1764399e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000001110100000101101010101111;
		b = 32'b01101111111111010001001110101011;
		correct = 32'b00110010010011011111100110100001;
		#400 //7.653726e-38 * 1.5664697e+29 = 1.19893295e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110010101111011100111111001110;
		b = 32'b00111101101011101100110000011010;
		correct = 32'b00110001000000011001101010010011;
		#400 //2.2096994e-08 * 0.08535023 = 1.8859836e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010111010110011111110100011001;
		b = 32'b10001110011001110001111101111110;
		correct = 32'b10100110010001001100111000110010;
		#400 //239681070000000.0 * -2.8488111e-30 = -6.8280607e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101110101110001101101111110100;
		b = 32'b00011000101111110011001100011110;
		correct = 32'b00001000000010100001000100000101;
		#400 //8.406423e-11 * 4.9423958e-24 = 4.154787e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001001001001101000001111101101;
		b = 32'b01100110110111001100100010101011;
		correct = 32'b00110000100011111001101111100110;
		#400 //2.0043554e-33 * 5.2131115e+23 = 1.0448928e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010011110011010011001000101;
		b = 32'b11010010000010011011001000011000;
		correct = 32'b01001101000001100100011110101000;
		#400 //-0.0009523372 * -147849610000.0 = 140802690.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000011111110100110001010111010;
		b = 32'b01010010100101011101111000111101;
		correct = 32'b10010111000100101001010011010100;
		#400 //-1.4716346e-36 * 321839330000.0 = -4.736299e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100110101010101101111010101010;
		b = 32'b00011011101011101100001011000111;
		correct = 32'b11000010111010010100101010110010;
		#400 //-4.0345486e+23 * 2.8911757e-22 = -116.64589
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000111010111110111100100001111;
		b = 32'b01011011010001100101111100101011;
		correct = 32'b10100011001011010010101010110101;
		#400 //-1.6812231e-34 * 5.5836684e+16 = -9.387392e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010000001110111001010111011110;
		b = 32'b00111010110011010000100101100101;
		correct = 32'b00001011100101100011110111100101;
		#400 //3.69947e-29 * 0.0015643059 = 5.7871027e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101011110010010111111010010100;
		b = 32'b10110110101010101010000111111010;
		correct = 32'b01100011000001100100110110001100;
		#400 //-4.8718368e+26 * -5.0852514e-06 = 2.4774515e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011110001101101110011111010100;
		b = 32'b11000000100111101001000001111010;
		correct = 32'b01011111011000101001010010011101;
		#400 //-3.294934e+18 * -4.9551363 = 1.6326847e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111100101000001010011100011011;
		b = 32'b10001010010101100010111010101000;
		correct = 32'b01000111100001100110100011111000;
		#400 //-6.6732544e+36 * -1.03125e-32 = 68817.94
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100001011101010001000000000111;
		b = 32'b11101011111110011101010101101111;
		correct = 32'b01001101111011110010100011100111;
		#400 //-8.303044e-19 * -6.0406088e+26 = 501554400.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000101111101110011110001101100;
		b = 32'b01110001010001010101000001101110;
		correct = 32'b10110111101111101000111100101100;
		#400 //-2.3249964e-35 * 9.770525e+29 = -2.2716435e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101010011110101101111101000110;
		b = 32'b00111011010011110111000001000011;
		correct = 32'b01100110010010110100100010001101;
		#400 //7.582146e+25 * 0.0031652607 = 2.3999468e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110100101110100010111001011101;
		b = 32'b10011110001010010100101111011101;
		correct = 32'b00010011011101100011111110001111;
		#400 //-3.4678934e-07 * -8.962474e-21 = 3.1080902e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011100010110111001010101000000;
		b = 32'b11010110111000001100001011000010;
		correct = 32'b01110011110000001100100110100110;
		#400 //-2.4722849e+17 * -123563540000000.0 = 3.0548429e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111110101010101010111000101010;
		b = 32'b10111010011111110000110110101000;
		correct = 32'b00111001101010100000110010010111;
		#400 //-0.33336002 * -0.0009729513 = 0.00032434307
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101001001011010000000011000010;
		b = 32'b11000001111110110001110110110001;
		correct = 32'b11101011101010011011001111001111;
		#400 //1.3071734e+25 * -31.389498 = -4.1031517e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011111001000011101101110101101;
		b = 32'b00110000110100110000111010000101;
		correct = 32'b11010000100001010111000100111110;
		#400 //-1.1663106e+19 * 1.5356397e-09 = -17910330000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010011011011011000111000111110;
		b = 32'b11000111100101011111011110111101;
		correct = 32'b10011011100010110010100110101110;
		#400 //2.9983736e-27 * -76783.48 = -2.3022556e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111011011100010010110111111;
		b = 32'b10010101100110100110011101011010;
		correct = 32'b10011101100011111010001011011010;
		#400 //60965.746 * -6.2363165e-26 = -3.802017e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001000001100111011101000110110;
		b = 32'b01001100001101111011111101110000;
		correct = 32'b01010101000000010000000010000011;
		#400 //184040.84 * 48168384.0 = 8864950000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100000100110111100011010101000;
		b = 32'b01100101010001010001110011101001;
		correct = 32'b01000110011011111110001011101110;
		#400 //2.638948e-19 * 5.817747e+22 = 15352.732
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110001011101111010111101111011;
		b = 32'b10101000110010000010111001101110;
		correct = 32'b11011010110000011010111000000100;
		#400 //1.22647904e+30 * -2.2224596e-14 = -2.7258001e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011110001000011101100111110010;
		b = 32'b00110010000000110111100000011100;
		correct = 32'b10010000101001100011110011101101;
		#400 //-8.568339e-21 * 7.652513e-09 = -6.5569326e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110001111001000111100001010011;
		b = 32'b00010100101101010001011001001101;
		correct = 32'b11000111001000011001110011111010;
		#400 //-2.2626574e+30 * 1.8285126e-26 = -41372.977
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000100001101011000111000001;
		b = 32'b01110001011100000100010001000001;
		correct = 32'b11100010011111001101010100011101;
		#400 //-9.800304e-10 * 1.18974266e+30 = -1.165984e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101010000010111110100101101000;
		b = 32'b10100111010001100001011011101101;
		correct = 32'b01010001110110001000011000011100;
		#400 //-4.228573e+25 * -2.7490448e-15 = 116245365000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000010110010011100111111110100;
		b = 32'b00000001010000110010111001111011;
		correct = 32'b00000100100110011101111000001011;
		#400 //100.90616 * 3.5849192e-38 = 3.617404e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001000100010110101011110011111;
		b = 32'b10000001101110000111010000011100;
		correct = 32'b10001010110010001100110001011010;
		#400 //285372.97 * -6.7757534e-38 = -1.9336168e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100010101111101110101100110100;
		b = 32'b10111101100001011101000011011010;
		correct = 32'b00100000110001111001011111100111;
		#400 //-5.1748634e-18 * -0.06533976 = 3.3812432e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100111011000011111000000001110;
		b = 32'b10101010010110100000010111111001;
		correct = 32'b10010010010000000110101110110001;
		#400 //3.1355156e-15 * -1.9364362e-13 = -6.0717257e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100010110001101101101011010010;
		b = 32'b10010111000101000110110111011010;
		correct = 32'b10111010011001101001011110101100;
		#400 //1.8341115e+21 * -4.796003e-25 = -0.00087964046
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000111011110000100101110100011;
		b = 32'b10111101100110011001001011100100;
		correct = 32'b10000101100101001111001110101101;
		#400 //1.8679674e-34 * -0.0749872 = -1.4007365e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011001110100101100100111111;
		b = 32'b10110011110101100001100110111010;
		correct = 32'b00111111100110111101100101010101;
		#400 //-12212543.0 * -9.969831e-08 = 1.21757
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011110011000110010111001001000;
		b = 32'b10101111000001000101011000100010;
		correct = 32'b11001101111010101110000010011010;
		#400 //4.0925252e+18 * -1.203593e-10 = -492573500.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111110001101101001010011010100;
		b = 32'b00101000010000000111110100110111;
		correct = 32'b10100111000010010100100011101101;
		#400 //-0.17830211 * 1.0685293e-14 = -1.9052102e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010111100001100101000010000111;
		b = 32'b10110011001110101100001111000100;
		correct = 32'b10001011010000111111101001110001;
		#400 //8.679875e-25 * -4.3484548e-08 = -3.7744045e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000110101010101111011011100010;
		b = 32'b00000111011000111101000101111100;
		correct = 32'b00001110100110000010010011010001;
		#400 //21883.441 * 1.7139144e-34 = 3.7506346e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000101101100001011101011010111;
		b = 32'b00000100101101110111000110111111;
		correct = 32'b10001010111111010100100000101100;
		#400 //-5655.355 * 4.3127553e-36 = -2.4390162e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001110010110011100011110001000;
		b = 32'b01101110100101010110001110101100;
		correct = 32'b00111101011111100010101111011001;
		#400 //2.6843386e-30 * 2.3116881e+28 = 0.062053535
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110011000011110011100100101111;
		b = 32'b01100000001001000000101001011101;
		correct = 32'b11010011101101111000110011011101;
		#400 //-3.334679e-08 * 4.728145e+19 = -1576684600000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011011100010101111101001000111;
		b = 32'b11011101011011001101101011001011;
		correct = 32'b01111001100000001001010110000001;
		#400 //-7.823746e+16 * -1.06669856e+18 = 8.345579e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101010000101110111110101100100;
		b = 32'b10111010010000011101000101011101;
		correct = 32'b01100100111001010110001011011010;
		#400 //-4.5784985e+25 * -0.0007393563 = 3.385142e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001000010111100111100000101001;
		b = 32'b10010010110000100111010001000110;
		correct = 32'b00011011101010001111110000011010;
		#400 //-227808.64 * -1.2271785e-27 = 2.7956185e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111100000010010001111001011110;
		b = 32'b00111010111011111011011000000101;
		correct = 32'b00110111100000000110010011011000;
		#400 //0.0083690565 * 0.0018288499 = 1.5305748e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111001001010001100000101001111;
		b = 32'b10111110000111011111110001101101;
		correct = 32'b01110111110100000100100111100111;
		#400 //-5.4764165e+34 * -0.15428324 = 8.4491927e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111010111001001000010011001110;
		b = 32'b00010100010000101111001001011110;
		correct = 32'b01001111101011100000010011111110;
		#400 //5.9326864e+35 * 9.8422955e-27 = 5839125500.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000110011100100010100111000;
		b = 32'b10101010110001001110101010100110;
		correct = 32'b00011100000111101010101000010000;
		#400 //-1.5008146e-09 * -3.4979414e-13 = 5.2497615e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100110000100001111001100001011;
		b = 32'b11000111111110111110001111000011;
		correct = 32'b11101110100011101001111101000010;
		#400 //1.7112603e+23 * -128967.52 = -2.20697e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110001100101101010110011011101;
		b = 32'b00100011100011010011011010001010;
		correct = 32'b10010101101001100011101010011111;
		#400 //-4.385227e-09 * 1.5310349e-17 = -6.7139354e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010010111001011101011100101100;
		b = 32'b00001011110110101101011111000000;
		correct = 32'b10011111010001000111101011110000;
		#400 //-493578750000.0 * 8.429517e-32 = -4.1606306e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101011100111101000011000000001;
		b = 32'b10001000101111011001110000111100;
		correct = 32'b00110100111010101101001101011011;
		#400 //-3.832862e+26 * -1.1411754e-33 = 4.3739678e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011110001110011111000000110101;
		b = 32'b01000111110000100001101110000011;
		correct = 32'b10100110100011001111110000000100;
		#400 //-9.843492e-21 * 99383.02 = -9.78276e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111100000101001001101000001111;
		b = 32'b11011001100101100001110111101100;
		correct = 32'b01010110001011100100011101000110;
		#400 //-0.009069934 * -5281768000000000.0 = 47905285000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001110111101100100011101111111;
		b = 32'b00110010111110010010011000001000;
		correct = 32'b00000010011011111011000000100001;
		#400 //6.071253e-30 * 2.900471e-08 = 1.7609493e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101111110011000110011111100101;
		b = 32'b10111001000110100000010101111001;
		correct = 32'b10101001011101011111010110111101;
		#400 //3.7181205e-10 * -0.00014688623 = -5.4614072e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111001111110001110011000110101;
		b = 32'b00011100011110011111010010010110;
		correct = 32'b01010110111100110000010110110111;
		#400 //1.6154485e+35 * 8.270331e-22 = 133602935000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111011101100011110110001010011;
		b = 32'b11100011100111100001010100100100;
		correct = 32'b11011111110110111011110100011001;
		#400 //0.0054297834 * -5.832218e+21 = -3.1667679e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000001111001000011101010100011;
		b = 32'b01000110111101011000101101000000;
		correct = 32'b10001001010110101110100001000011;
		#400 //-8.383811e-38 * 31429.625 = -2.6350004e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100100100111011000000101111011;
		b = 32'b10011000010110101100001011001001;
		correct = 32'b10111101100001101001100000011011;
		#400 //2.324375e+22 * -2.8274181e-24 = -0.065719806
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110001010011001001001111010;
		b = 32'b11100111101100100010011011101011;
		correct = 32'b01011110011011000000001101000000;
		#400 //-2.5268223e-06 * -1.6825983e+24 = 4.2516267e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001101010001010010111110110010;
		b = 32'b00111011100000001011011101011101;
		correct = 32'b01001001010001100100101000101011;
		#400 //206764830.0 * 0.0039281086 = 812194.7
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101110010001100111011101111000;
		b = 32'b10001011000101001010101111101111;
		correct = 32'b10111001111001101000010010111001;
		#400 //1.5355615e+28 * -2.8633112e-32 = -0.00043967905
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001001010100010000010011111100;
		b = 32'b00100100010111100110110101010100;
		correct = 32'b10101110001101011001101110010110;
		#400 //-856143.75 * 4.823118e-17 = -4.1292823e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110011111001111011110011111100;
		b = 32'b01100101100100001010101100001010;
		correct = 32'b01011010000000101111010100100010;
		#400 //1.0791152e-07 * 8.539699e+22 = 9215318000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100001000100011001001001011111;
		b = 32'b11101101001101010010011111000110;
		correct = 32'b11001110110011100000011000110110;
		#400 //4.932163e-19 * -3.5040544e+27 = -1728256800.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000100101110100100010001111000;
		b = 32'b01010011001101011101111011100100;
		correct = 32'b00011000100001000101010010010110;
		#400 //4.379127e-36 * 781128560000.0 = 3.420661e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110100010001010000000100110100;
		b = 32'b01000010000010101010011110010100;
		correct = 32'b11110110110101010110011100110111;
		#400 //-6.243328e+31 * 34.66365 = -2.1641654e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100111000100101101000011000110;
		b = 32'b00111110011111101000011010110111;
		correct = 32'b01100110000100011111100001100111;
		#400 //6.933167e+23 * 0.24856077 = 1.7233134e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111000101100000111000001101001;
		b = 32'b10100001001101001001010010111010;
		correct = 32'b01011010011110001110101100010110;
		#400 //-2.862888e+34 * -6.118321e-19 = 1.7516068e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001010000111011101010001101111;
		b = 32'b00101011011111111111101011010000;
		correct = 32'b00110110000111011101000100111100;
		#400 //2585883.8 * 9.094227e-13 = 2.3516614e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000110000000111101111110001001;
		b = 32'b01100100011100100011001110001111;
		correct = 32'b11101010111110011000011110111101;
		#400 //-8439.884 * 1.7871309e+22 = -1.5083177e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111011100111000000011100101000;
		b = 32'b00101110010011101100111000000110;
		correct = 32'b11101010011111000001011010100111;
		#400 //-1.6202869e+36 * 4.7021963e-11 = -7.618907e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100111000000101011011010011100;
		b = 32'b10111110110001011001100010010001;
		correct = 32'b11100110010010011100100011011001;
		#400 //6.172762e+23 * -0.3859296 = -2.3822516e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110011011101110101101101010101;
		b = 32'b10000011000010011100101001111100;
		correct = 32'b10110111000001010010001110000110;
		#400 //1.9597622e+31 * -4.049312e-37 = -7.935689e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011100011111111011101100000111;
		b = 32'b01011010110000001110110001101010;
		correct = 32'b00110111110000001011100001110000;
		#400 //8.461415e-22 * 2.7151568e+16 = 2.2974069e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110101100001000001000000101010;
		b = 32'b00000001010111101000111100111100;
		correct = 32'b00110111011001011001111111010001;
		#400 //3.3481984e+32 * 4.0877726e-38 = 1.3686674e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010000101111011010101000110011;
		b = 32'b11101100110011000011010010011111;
		correct = 32'b00111110000101110100101010011101;
		#400 //-7.480959e-29 * -1.9749549e+27 = 0.14774556
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101110111001001111011000011010;
		b = 32'b10011001111000111101000101101110;
		correct = 32'b01001001010010111100000110001000;
		#400 //-3.543005e+28 * -2.3555838e-23 = 834584.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011111011110001110011001010010;
		b = 32'b01100110101001011010110101001001;
		correct = 32'b01000110101000010001010011101101;
		#400 //5.270656e-20 * 3.911935e+23 = 20618.463
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011000001000101011011011110111;
		b = 32'b00011110111010010001001011100101;
		correct = 32'b00110111100101000010010010001001;
		#400 //715626850000000.0 * 2.4677649e-20 = 1.7659988e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100110111101010110111100011010;
		b = 32'b10101001000100011100101101011001;
		correct = 32'b10010000100010111100011011100010;
		#400 //1.7030404e-15 * -3.2372844e-14 = -5.513226e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010011001100100001110110100011;
		b = 32'b11101010111110111100101101111001;
		correct = 32'b01111110101011110011000010100001;
		#400 //-765001400000.0 * -1.5220063e+26 = 1.164337e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101110101011100001100001100111;
		b = 32'b11011101111010101010011010011011;
		correct = 32'b01001101000111111001001110011011;
		#400 //-7.9169386e-11 * -2.1135465e+18 = 167328180.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111011110011101100010010001;
		b = 32'b10001011010010101100100100110010;
		correct = 32'b00000011010001011110100100111110;
		#400 //-1.489198e-05 * -3.9055147e-32 = 5.8160846e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100000111011111100101101000111;
		b = 32'b10000110110011101110110010001010;
		correct = 32'b00101000010000011101001100100100;
		#400 //-1.3823186e+20 * -7.783615e-35 = 1.0759436e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100100011011100011110110110110;
		b = 32'b00111001011000001010000111001010;
		correct = 32'b10011110010100010000110010010000;
		#400 //-5.1660295e-17 * 0.00021422576 = -1.1066966e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010111010100010011110101100011;
		b = 32'b10010000110010101010100101010000;
		correct = 32'b10101000101001011010010011010011;
		#400 //230061580000000.0 * -7.993582e-29 = -1.8390161e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111100010011000111101110010111;
		b = 32'b01111011001011001011001011110111;
		correct = 32'b11111000000010011111000111111101;
		#400 //-0.012480638 * 8.967049e+35 = -1.119145e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101111001011101011011111111000;
		b = 32'b00100011000010011011110001010101;
		correct = 32'b00010010101111000000000111111010;
		#400 //1.5890567e-10 * 7.466666e-18 = 1.1864955e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101001111111011111110001000101;
		b = 32'b01001101100100110010101000011110;
		correct = 32'b01111000000100100000000110100101;
		#400 //3.8381193e+25 * 308626370.0 = 1.1845448e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000011111110001001101011011011;
		b = 32'b10000001100111010000110000000011;
		correct = 32'b00000110000110001000001010100010;
		#400 //-497.2098 * -5.768993e-38 = 2.8683996e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100001001011110100010000000010;
		b = 32'b10001111110100010001000001100000;
		correct = 32'b10110001100011110010000110111100;
		#400 //2.0206754e+20 * -2.0615299e-29 = -4.165683e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101000000011101100111001110110;
		b = 32'b00100111001110101000100010100010;
		correct = 32'b00001111110100000001110001110100;
		#400 //7.9273526e-15 * 2.5886754e-15 = 2.0521343e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101010111110011000010010001101;
		b = 32'b00001100111001000100011101000111;
		correct = 32'b00111000010111100111111110000111;
		#400 //1.5082424e+26 * 3.517186e-31 = 5.3047694e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001000011010111110001101100111;
		b = 32'b00010010110001111011000001110101;
		correct = 32'b10011011101110000000000001011101;
		#400 //-241549.61 * 1.2602166e-27 = -3.0440481e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010101111010111011010101000111;
		b = 32'b10100100011010001100000100000111;
		correct = 32'b10111010110101100100111000000010;
		#400 //32395477000000.0 * -5.047048e-17 = -0.0016350152
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010101110100110111110110011011;
		b = 32'b00110011010110101100000111100111;
		correct = 32'b00001001101101001011100100100111;
		#400 //8.542039e-26 * 5.0933433e-08 = 4.350754e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001011010000000111111010110010;
		b = 32'b11101110101010000010011000101111;
		correct = 32'b00111010011111001101111110110110;
		#400 //-3.707317e-32 * -2.6019821e+28 = 0.00096463726
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101010010000000001011100011101;
		b = 32'b10110000000110101000100000110000;
		correct = 32'b01011010111001111110100000101111;
		#400 //-5.8055727e+25 * -5.621841e-10 = 3.2638004e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101000111101101001101101011000;
		b = 32'b10001000011000110111111010101110;
		correct = 32'b00110001110110110010010111000111;
		#400 //-9.316542e+24 * -6.845924e-34 = 6.3780337e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000010000010011110110111101000;
		b = 32'b11011001100001000010101011110000;
		correct = 32'b00011100000011100110101110011100;
		#400 //-1.0133446e-37 * -4650238400000000.0 = 4.712294e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010010101101111100101011001000;
		b = 32'b11100000011110011101001101010001;
		correct = 32'b10110011101100110101101111110011;
		#400 //1.1598913e-27 * -7.2007285e+19 = -8.3520625e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011001000100010110011000011010;
		b = 32'b00111100001111110010011111011111;
		correct = 32'b01010101110110010010001110100101;
		#400 //2557883300000000.0 * 0.011667221 = 29843390000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100101000000100000010011001010;
		b = 32'b10101110011101101101101010000001;
		correct = 32'b11010011111110101011111100100111;
		#400 //3.837475e+22 * -5.6127995e-11 = -2153897700000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011011100111000001100111100101;
		b = 32'b10111111010001101100101001011110;
		correct = 32'b00011011011100100110111011011010;
		#400 //-2.582477e-22 * -0.7765254 = 2.0053589e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111111101111110000100101110100;
		b = 32'b01101111101000111101010001000100;
		correct = 32'b01101111111101001000001011010111;
		#400 //1.492476 * 1.0140534e+29 = 1.5134504e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010011101010110001011101001101;
		b = 32'b11001000100100111110011000011011;
		correct = 32'b00011100110001011011000001010100;
		#400 //-4.3189445e-27 * -302896.84 = 1.3081946e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011111000111010001011000001;
		b = 32'b00100110101111010100110101011001;
		correct = 32'b10110011001010000101001111110000;
		#400 //-29836674.0 * 1.3135475e-15 = -3.919189e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001010111010110111101100000100;
		b = 32'b01011000110110010101101000000011;
		correct = 32'b11100100010001111110111000010010;
		#400 //-7716226.0 * 1911845000000000.0 = -1.4752227e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011010000100101100000001011011;
		b = 32'b01010100100100100000001001011010;
		correct = 32'b11101111001001110110011000011010;
		#400 //-1.0326711e+16 * 5016837400000.0 = -5.180743e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110011100000111101110011001001;
		b = 32'b01111000101001010110010001000101;
		correct = 32'b01101100101010100110000111100111;
		#400 //6.1403234e-08 * 2.6836334e+34 = 1.6478378e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110100100011010010101001110001;
		b = 32'b10010001010011001101111000110110;
		correct = 32'b11000110011000011111000010110101;
		#400 //8.947445e+31 * -1.6161236e-28 = -14460.177
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011001110101100011111000111011;
		b = 32'b00101111000011001010110010011101;
		correct = 32'b00001001011010110111010011111011;
		#400 //2.2152216e-23 * 1.279425e-10 = 2.83421e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111000011111100001101010011111;
		b = 32'b10100101010001010111110101100111;
		correct = 32'b10011110010001000000011011110110;
		#400 //6.0583112e-05 * -1.7129514e-16 = -1.0377593e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101000111010000101111111000111;
		b = 32'b01110100100000100111001110001100;
		correct = 32'b11011101111011001101001100001010;
		#400 //-2.5798711e-14 * 8.268337e+31 = -2.1331243e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000100111010110110001101000010;
		b = 32'b01010001111100110011111011110000;
		correct = 32'b00010111010111111010100100010110;
		#400 //5.533939e-36 * 130591620000.0 = 7.2268603e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000101000111111010111110011110;
		b = 32'b10001110101101111110011011101011;
		correct = 32'b00010100011001010110110100101001;
		#400 //-2554.976 * -4.533535e-30 = 1.15830735e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100110010110011010100000111010;
		b = 32'b11001000100001110000010101011111;
		correct = 32'b01101111011001011001100010001111;
		#400 //-2.5696419e+23 * -276522.97 = 7.10565e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011110000001110010000110111010;
		b = 32'b01000101100110100100101111011111;
		correct = 32'b01100100001000101110010010101101;
		#400 //2.434317e+18 * 4937.484 = 1.2019401e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001001100100011100100011111111;
		b = 32'b00100100111101001111111000110010;
		correct = 32'b10101111000010111000010001010101;
		#400 //-1194271.9 * 1.06248756e-16 = -1.268899e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111101101111000010010111110111;
		b = 32'b11010011000101101100111111110100;
		correct = 32'b11010001010111011010111000101010;
		#400 //0.09186929 * -647734000000.0 = -59506860000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010111011001110100101000100011;
		b = 32'b01010101001110111101011000101101;
		correct = 32'b01101101001010011011010010101000;
		#400 //254305600000000.0 * 12908035000000.0 = 3.2825854e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010101101101101000101111111000;
		b = 32'b11010101011001111101011000001000;
		correct = 32'b00101011101001010101000011101011;
		#400 //-7.3730046e-26 * -15931653000000.0 = 1.1746414e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010101101011011100001110011101;
		b = 32'b10011001000010011101011101010011;
		correct = 32'b00101111001110110001111110101101;
		#400 //-23881958000000.0 * -7.126218e-24 = 1.7018804e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110011100110001110111011010101;
		b = 32'b00000101100111110100010111101000;
		correct = 32'b10111001101111100100110000110011;
		#400 //-2.4233191e+31 * 1.4977968e-35 = -0.00036296397
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111000110100101111011010010110;
		b = 32'b01001001100101110111010000111110;
		correct = 32'b01000010111110011001111001111011;
		#400 //0.000100595105 * 1240711.8 = 124.80953
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010111011010111001010101010;
		b = 32'b10101100100101101100100110011011;
		correct = 32'b00101000000010111101110000101110;
		#400 //-0.0018115838 * -4.285639e-12 = 7.763794e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111111011011111011101110001101;
		b = 32'b00011000001111011100100010010111;
		correct = 32'b01011000001100011011100101001111;
		#400 //3.1865931e+38 * 2.452895e-24 = 781637800000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110101001100110000011001010111;
		b = 32'b10001111010100000110110110110011;
		correct = 32'b01000101000100011100000111011110;
		#400 //-2.2694085e+32 * -1.0276319e-29 = 2332.1167
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011000000011000100001110011101;
		b = 32'b11100101000111001100110111011110;
		correct = 32'b00111101101010111101001111111111;
		#400 //-1.8128712e-24 * -4.628042e+22 = 0.083900444
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000100111011100111101001100111;
		b = 32'b01001011101010101010100101000011;
		correct = 32'b10010001000111101111101011110110;
		#400 //-5.606594e-36 * 22368902.0 = -1.2541336e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010010100000100100001010100111;
		b = 32'b01111000101000010000010100110100;
		correct = 32'b01001011101000111101110100100010;
		#400 //8.2205845e-28 * 2.6127041e+34 = 21477956.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111110011111011000101101111111;
		b = 32'b10101101111001010101001111011111;
		correct = 32'b11101100111000110010000011011010;
		#400 //8.4254747e+37 * -2.6071532e-11 = -2.1966504e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010101110111111000100110010111;
		b = 32'b11111011011000101011001101101101;
		correct = 32'b11010001110001011111010000100100;
		#400 //9.028606e-26 * -1.1770983e+36 = -106275570000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110110011011001010100000010111;
		b = 32'b01101010010001011011100010111100;
		correct = 32'b01100001001101101100100000100000;
		#400 //3.5264582e-06 * 5.9757692e+25 = 2.10733e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001110011010100111001111100010;
		b = 32'b11001011110000101010000001010110;
		correct = 32'b11011010101100100011111010101000;
		#400 //983365760.0 * -25510060.0 = -2.5085719e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101101111111001011010010000111;
		b = 32'b10001100100111011001011001100001;
		correct = 32'b00111011000110111000111100101000;
		#400 //-9.7760583e+27 * -2.4280186e-31 = 0.002373645
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001001100011000000101001000011;
		b = 32'b10110110010101000101011110001011;
		correct = 32'b01000000011010000101000011000110;
		#400 //-1147208.4 * -3.1641418e-06 = 3.62993
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111100011101011100110010100100;
		b = 32'b10011000011001110110100010001110;
		correct = 32'b00010101010111100011000000001011;
		#400 //-0.015002403 * -2.9908837e-24 = 4.4870442e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000110011111111110100101001111;
		b = 32'b00111100101001000100100111101011;
		correct = 32'b10000011101001000011101101011011;
		#400 //-4.8131578e-35 * 0.020054778 = -9.652681e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101000111011000010111100101100;
		b = 32'b00101011011011110011101011100000;
		correct = 32'b10010100110111001011011001011011;
		#400 //-2.6221721e-14 * 8.499156e-13 = -2.228625e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111100010011110001011100111100;
		b = 32'b10011101101000010111000111010110;
		correct = 32'b01011010100000101001100110110011;
		#400 //-4.3011068e+36 * -4.273405e-21 = 1.838037e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100111100010101101001000110111;
		b = 32'b00100000000111100100001100110010;
		correct = 32'b01001000001010111010010001011100;
		#400 //1.3111287e+24 * 1.3405354e-19 = 175761.44
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110101110011000000100010011010;
		b = 32'b10011100010100010110111011100001;
		correct = 32'b01010010101001101110101101100101;
		#400 //-5.1728663e+32 * -6.9295607e-22 = 358456920000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001010000101001011010010001001;
		b = 32'b10011100000010011010110000110110;
		correct = 32'b10100110100111111111000101001100;
		#400 //2436386.2 * -4.5552075e-22 = -1.1098245e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001001111101100111101101011100;
		b = 32'b00011011110001001101000011010011;
		correct = 32'b00100110001111010111111110000010;
		#400 //2019179.5 * 3.256043e-22 = 6.5745353e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001010111010100100100011001011;
		b = 32'b10111001001010111101111110111011;
		correct = 32'b10000100100111010100101101100000;
		#400 //2.2560762e-32 * -0.00016391177 = -3.6979744e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010001101011101101101011010001;
		b = 32'b10001000010100100010101001101100;
		correct = 32'b00011010100011111000110001111001;
		#400 //-93874430000.0 * -6.3244443e-34 = 5.937036e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110101000111010010110000010111;
		b = 32'b10100010001000010000101011000000;
		correct = 32'b01010111110001011011111010101000;
		#400 //-1.9923947e+32 * -2.182526e-18 = 434845300000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001110110111010111110111101000;
		b = 32'b10010100010111000010110010010101;
		correct = 32'b00100011101111100111111011000110;
		#400 //-1858008000.0 * -1.1115954e-26 = 2.0653532e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000101101100110011101100001011;
		b = 32'b01111011101111011100101000110110;
		correct = 32'b11000010000001001110000000101010;
		#400 //-1.6854768e-35 * 1.9708909e+36 = -33.21891
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101010100101010010111111001010;
		b = 32'b00011110111101011011011001001011;
		correct = 32'b01001010000011110011000011111000;
		#400 //9.017781e+25 * 2.6015779e-20 = 2346046.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111000110010100111011000000001;
		b = 32'b11000001011110001011111101010010;
		correct = 32'b11111010110001001011100110100000;
		#400 //3.2851168e+34 * -15.546709 = -5.1072755e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110000001010101010100100010000;
		b = 32'b10011111101100100000110100001110;
		correct = 32'b10010000011011010110010010000010;
		#400 //6.208589e-10 * -7.540753e-20 = -4.6817437e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101110110100110111010010000000;
		b = 32'b11000001000100001011011100011001;
		correct = 32'b01110000011011110001000110001010;
		#400 //-3.2721088e+28 * -9.044702 = 2.9595248e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101011110100011101011101011101;
		b = 32'b10010100010101011101110100111010;
		correct = 32'b00000000101011110100110110000111;
		#400 //-1.4910118e-12 * -1.0797381e-26 = 1.6099023e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111111110010000111000001110011;
		b = 32'b11010001111001010101010001011101;
		correct = 32'b11010010001100111000111010100101;
		#400 //1.5659317 * -123120360000.0 = -192798080000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100011100101001000010001100001;
		b = 32'b00011101011111100001111000101001;
		correct = 32'b10000001100100110110110011011000;
		#400 //-1.6102257e-17 * 3.3632213e-21 = -5.4155455e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111101001110001100010101010001;
		b = 32'b00101001111100001100111100111011;
		correct = 32'b10100111101011011100111010001110;
		#400 //-0.04511005 * 1.069409e-13 = -4.8241093e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100000100111111111011001000111;
		b = 32'b01111101001111110010000001000100;
		correct = 32'b11011110011011101101100111010000;
		#400 //-2.709862e-19 * 1.587813e+37 = -4.302754e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011001011110011111000001011001;
		b = 32'b01001110111110010100011100110110;
		correct = 32'b10101000111100110110000001001101;
		#400 //-1.2921536e-23 * 2091096800.0 = -2.7020183e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101010001001100000110111100011;
		b = 32'b00011010100010001010110111010101;
		correct = 32'b11000101001100010101000001000100;
		#400 //-5.0186816e+25 * 5.652912e-23 = -2837.0166
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010101010111000000001111011101;
		b = 32'b11000110111111110100100010100100;
		correct = 32'b10011100110110110110011001000111;
		#400 //4.4431694e-26 * -32676.32 = -1.4518642e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110011000110000100000110001;
		b = 32'b01101001110011011000000000001010;
		correct = 32'b11100000101101100011111100011100;
		#400 //-3.3830404e-06 * 3.1054305e+25 = -1.0505797e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111111110100010011100110111011;
		b = 32'b00101110111000111110100010001000;
		correct = 32'b00101111001110100100010000111100;
		#400 //1.6345743 * 1.0364071e-10 = 1.6940843e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101010110001010010011101110010;
		b = 32'b10101110011000011001101111001110;
		correct = 32'b11011001101011011011111110101001;
		#400 //1.1917233e+26 * -5.129746e-11 = -6113238000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000011100010001110011001111111;
		b = 32'b01011101001101110101100111000001;
		correct = 32'b10100001010001000001100110001000;
		#400 //-8.046281e-37 * 8.257377e+17 = -6.6441173e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100100001111000110101010110111;
		b = 32'b11110000000010010010001100000000;
		correct = 32'b01010100110010011101110110111101;
		#400 //-4.0856393e-17 * -1.6976703e+29 = 6936068600000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110101011100101011001010111010;
		b = 32'b10010011000010011000111001100101;
		correct = 32'b00001001000000100110100010100100;
		#400 //-9.0412107e-07 * -1.7362037e-27 = 1.5697383e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111001110010101111011000110100;
		b = 32'b11011000101010001010101011110000;
		correct = 32'b11010011000001011011100100011000;
		#400 //0.00038711878 * -1483617000000000.0 = -574336000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000000000101000000001011111101;
		b = 32'b11111011111011000111111011101101;
		correct = 32'b10111011100100111110010101101010;
		#400 //1.837782e-39 * -2.4559128e+36 = -0.0045134323
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110100100010110111011101001100;
		b = 32'b00001111011100000001001111101010;
		correct = 32'b10000100100000101100101010110001;
		#400 //-2.5977567e-07 * 1.1836749e-29 = -3.0748996e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000001010110110011000101011100;
		b = 32'b10110011000011100101100101110011;
		correct = 32'b10110100111100111100001111101111;
		#400 //13.699551 * -3.3143305e-08 = -4.5404838e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100010101001100001000001000001;
		b = 32'b01010010110000100110011111100101;
		correct = 32'b11110101111111000011011101101101;
		#400 //-1.5316654e+21 * 417483360000.0 = -6.394448e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111100011110100001100010100111;
		b = 32'b00000001001011100001111001011010;
		correct = 32'b00111110001010100001101001101000;
		#400 //5.194297e+36 * 3.198053e-38 = 0.16611636
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001100001101101000001100110110;
		b = 32'b11001111011001110001000101000010;
		correct = 32'b11011100001001001011110010110011;
		#400 //47844570.0 * -3876668000.0 = -1.854775e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110111100111010000100100100100;
		b = 32'b00110001010111110110011011000110;
		correct = 32'b11101001100010010000101000000001;
		#400 //-6.370125e+33 * 3.250919e-09 = -2.070876e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101101110110110110000110110110;
		b = 32'b10001100011010100100101111110100;
		correct = 32'b10111010110010001100100001100111;
		#400 //8.486918e+27 * -1.8049561e-31 = -0.0015318514
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011010100001100100011110011;
		b = 32'b10001000110101100010001010101011;
		correct = 32'b00010100101011101010010001000001;
		#400 //-13682931.0 * -1.2887807e-33 = 1.7634297e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011010100110011001101110010001;
		b = 32'b10111001101010111111100101000011;
		correct = 32'b10010100110011100110000011110101;
		#400 //6.353065e-23 * -0.00032801376 = -2.0838927e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110101111111001001111010110100;
		b = 32'b11000100010001110011110100110011;
		correct = 32'b11111010110001001001101111000010;
		#400 //6.4046762e+32 * -796.95624 = -5.1042466e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000011010011001110111111110001;
		b = 32'b10110010000100110011001110010011;
		correct = 32'b10110101111010111010111000100010;
		#400 //204.93727 * -8.568253e-09 = -1.7559544e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110001010010011001100100001011;
		b = 32'b00111011001100111011111000111101;
		correct = 32'b10101101000011011000101111010010;
		#400 //-2.9336344e-09 * 0.0027426623 = -8.045968e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001111010001001100100011100111;
		b = 32'b01101011110001100011100110010010;
		correct = 32'b10111011100110000101111110100100;
		#400 //-9.7022385e-30 * 4.7927836e+26 = -0.004650073
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000101011000011000110011111001;
		b = 32'b01100110111011101000000011011000;
		correct = 32'b01101100110100100010001010010100;
		#400 //3608.8108 * 5.6315e+23 = 2.0323017e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110100000000011011000111100110;
		b = 32'b10111101110110110111001101011011;
		correct = 32'b11110010010111100101101101000010;
		#400 //4.110196e+31 * -0.10715362 = -4.4042238e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110110100011100111010111001101;
		b = 32'b10100111010000101101101110111001;
		correct = 32'b10011110010110001101111100010110;
		#400 //4.2456436e-06 * -2.704202e-15 = -1.1481078e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011000010000111001101100100001;
		b = 32'b00111010010010100110011111100100;
		correct = 32'b10010011000110101010011111001010;
		#400 //-2.528148e-24 * 0.00077211694 = -1.952026e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011110101011101000000000000;
		b = 32'b01000000110101101101000110010000;
		correct = 32'b11001101001100110110101011100111;
		#400 //-28024832.0 * 6.7130814 = -188132980.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011001010000011001111100111011;
		b = 32'b10110111001111110101101000110011;
		correct = 32'b01010001000100001011101000000110;
		#400 //-3406234100000000.0 * -1.1405488e-05 = 38849765000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011001101100100001001010000101;
		b = 32'b11101110111111111110101101010101;
		correct = 32'b01001001001100100000010000100101;
		#400 //-1.8412249e-23 * -3.9601588e+28 = 729154.3
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010010111000010000111011001011;
		b = 32'b10111110001000010000110001100101;
		correct = 32'b10010001100011011001010100110011;
		#400 //1.4203143e-27 * -0.15727384 = -2.2337829e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100011110100001000101111010110;
		b = 32'b00011101100001010111110111011001;
		correct = 32'b01000001110110010111111001010110;
		#400 //7.693998e+21 * 3.533493e-21 = 27.186687
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110100011111011110010010101101;
		b = 32'b11100001101010110110010100001001;
		correct = 32'b11010110101010011111101111110100;
		#400 //2.3645653e-07 * -3.952092e+20 = -93449800000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110100110000001011110000111001;
		b = 32'b00001111110010010001110000111100;
		correct = 32'b01000101000101110110100100001011;
		#400 //1.2216047e+32 * 1.9831006e-29 = 2422.5652
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010000100110011100110010101100;
		b = 32'b11100111001101000010110100100000;
		correct = 32'b11111000010110000111111000001010;
		#400 //20642620000.0 * -8.508584e+23 = -1.7563945e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010100111000110000101101101110;
		b = 32'b11100000100000011111100011001100;
		correct = 32'b10110101111001101000101011010101;
		#400 //2.292565e-26 * -7.492368e+19 = -1.7176741e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010000100001101011011010010111;
		b = 32'b11000110111101001110010011111100;
		correct = 32'b11011000000000001101111010000111;
		#400 //18080905000.0 * -31346.492 = -566772940000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110110010111111111101000101101;
		b = 32'b00001001110111100010110010000100;
		correct = 32'b00000000110000100110000111100110;
		#400 //3.337521e-06 * 5.348642e-33 = 1.7851206e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010110101110001000100100010100;
		b = 32'b01010010000101111000010101010100;
		correct = 32'b10101001010110100111000111101101;
		#400 //-2.9813312e-25 * 162694230000.0 = -4.850454e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011000000111110011101101011101;
		b = 32'b01100111110001101011110100100000;
		correct = 32'b11000000011101110011101100011001;
		#400 //-2.058024e-24 * 1.8770346e+24 = -3.862982
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110001010000011101101001101111;
		b = 32'b11111110110001000000011111001111;
		correct = 32'b11110000100101000111000100100111;
		#400 //2.8209362e-09 * -1.3028462e+38 = -3.675246e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001101011110110101010101001100;
		b = 32'b10111001110000111100100111111010;
		correct = 32'b10000111110000000011100001000100;
		#400 //7.744802e-31 * -0.00037343783 = -2.892202e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010001000001110010010101100011;
		b = 32'b10111101011011001100110100110101;
		correct = 32'b00001110111110100000010110011000;
		#400 //-1.0661143e-28 * -0.05781289 = 6.1635145e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110100010100111100011011001001;
		b = 32'b00100001111110000100110010111010;
		correct = 32'b11010110110011010110100000001100;
		#400 //-6.7114653e+31 * 1.6825443e-18 = -112923380000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111110110101111100100100000101;
		b = 32'b10110011000011110101110111100111;
		correct = 32'b01110010011100011011000011100001;
		#400 //-1.4341389e+38 * -3.3380186e-08 = 4.787182e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101101111001101110011101111000;
		b = 32'b00000011010100010000101111101110;
		correct = 32'b00110001101111001000110110111100;
		#400 //8.9326726e+27 * 6.1433274e-37 = 5.4876335e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111000111001010011101001101000;
		b = 32'b10110000110001100000000011111110;
		correct = 32'b01101010001100010100110000010000;
		#400 //-3.7194394e+34 * -1.4406678e-09 = 5.3584766e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001111110011010011000110001001;
		b = 32'b01010100110011000100101100000101;
		correct = 32'b00100101001000111011111110011011;
		#400 //2.0233641e-29 * 7019455600000.0 = 1.4202915e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101000011100001001101100111010;
		b = 32'b10011001111001101110001010000110;
		correct = 32'b00000010110110010000000001011101;
		#400 //-1.3356336e-14 * -2.3872935e-23 = 3.1885493e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000011010100001011000011111101;
		b = 32'b11110100101000110000110000101110;
		correct = 32'b00111000100001001110101010011111;
		#400 //-6.132888e-37 * -1.0334368e+32 = 6.337952e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010101011110001101011111010110;
		b = 32'b11000101100110011000111110100000;
		correct = 32'b01011011100101010100010010011011;
		#400 //-17100368000000.0 * -4913.953 = 8.403041e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101001000101011111101100011011;
		b = 32'b11011001010000000010001001100010;
		correct = 32'b11000010111000010010000011110010;
		#400 //3.3302445e-14 * -3380062500000000.0 = -112.56435
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011000101000101110001110011100;
		b = 32'b00101111101101111100011000111011;
		correct = 32'b10001000111010011101110110101100;
		#400 //-4.2105845e-24 * 3.3428357e-10 = -1.4075292e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100000100011000001000001010010;
		b = 32'b11101111001000111100001110111110;
		correct = 32'b01010000001100110011001011111001;
		#400 //-2.3727722e-19 * -5.0682694e+28 = 12025849000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100010000110000100011111001;
		b = 32'b01000111100101000101100101111001;
		correct = 32'b01001100011000100000101010110101;
		#400 //780.1402 * 75954.945 = 59255508.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111101011111001101011010100001;
		b = 32'b00101000111001001100010110000111;
		correct = 32'b11100110111000011111001000111110;
		#400 //-2.1004992e+37 * 2.5398749e-14 = -5.3350052e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111111110101010110001011101010;
		b = 32'b00001001010100000110010110000100;
		correct = 32'b00001001101011011011010011111100;
		#400 //1.6670811 * 2.5084822e-33 = 4.1818432e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100011011001000011010100011100;
		b = 32'b11010010001010000010010100111101;
		correct = 32'b00110110000101011110010000001100;
		#400 //-1.2371151e-17 * -180544820000.0 = 2.233547e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010111011011101111001101011101;
		b = 32'b01101100100111101011011010100101;
		correct = 32'b11000100100101000010010010101110;
		#400 //-7.7209115e-25 * 1.5349824e+27 = -1185.1462
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000111110111011110100101101;
		b = 32'b01110101101111101110100000101010;
		correct = 32'b11100111001110111011101010110100;
		#400 //-1.8316421e-09 * 4.8400647e+32 = -8.865266e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110001101111110111011011111000;
		b = 32'b01001001110011110100000100101001;
		correct = 32'b11111100000110110000000111101110;
		#400 //-1.8961748e+30 * 1697829.1 = -3.2193806e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011111100000101101110000110011;
		b = 32'b10100110101111010010111000001001;
		correct = 32'b00000110110000010110100000110100;
		#400 //-5.542143e-20 * -1.3126987e-15 = 7.2751644e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110111001101001110111111111;
		b = 32'b00001101100111100111100000111000;
		correct = 32'b10000101000011101100000111010000;
		#400 //-6.8729273e-06 * 9.766443e-31 = -6.712406e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000101111100111001100001000110;
		b = 32'b01100100011101011110011000001011;
		correct = 32'b00101010111010011111101110100000;
		#400 //2.2907547e-35 * 1.8144115e+22 = 4.1563714e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111111111110110100101010000110;
		b = 32'b00000110010011110000110100010110;
		correct = 32'b01111111111110110100101010000110;
		#400 //nan * 3.8941987e-35 = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011010001110110110101111001000;
		b = 32'b00111010011011000101101111100110;
		correct = 32'b10010101001011010000101010100100;
		#400 //-3.875776e-23 * 0.00090163795 = -3.4945466e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010100000100001001101001111000;
		b = 32'b10101101100011011101000011001000;
		correct = 32'b00000010001000000011011000000101;
		#400 //-7.300606e-27 * -1.6122562e-11 = 1.1770446e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101010000001110110101110001010;
		b = 32'b00000001001011010001001100110001;
		correct = 32'b00101011101101110001101110100110;
		#400 //4.0928206e+25 * 3.178885e-38 = 1.3010606e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101011100100000010111100100101;
		b = 32'b11100000111000111110001000101100;
		correct = 32'b11001101000000000101100100110000;
		#400 //1.0244901e-12 * -1.31365885e+20 = -134583040.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110011100101101110001101011000;
		b = 32'b00100000110010110011011111000011;
		correct = 32'b11010100111011111000111001001001;
		#400 //-2.3909168e+31 * 3.4426438e-19 = -8231074700000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000110111001111100101110101101;
		b = 32'b01101011001100100110000000101111;
		correct = 32'b00110010101000011000001010110101;
		#400 //8.7191817e-35 * 2.1564301e+26 = 1.8802305e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111011010011100010100001011011;
		b = 32'b00001010010101111011011011101000;
		correct = 32'b01000110001011011011011100110000;
		#400 //1.07043166e+36 * 1.0386274e-32 = 11117.797
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100011111100000100110110101111;
		b = 32'b01110110000011001100111001000110;
		correct = 32'b11011010100001000010110000011100;
		#400 //-2.6053752e-17 * 7.1397e+32 = -1.8601598e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011110010100110001000011111001;
		b = 32'b00110101110100101101100111000000;
		correct = 32'b11010100101011011101011101110100;
		#400 //-3.8022324e+18 * 1.5709593e-06 = -5973152400000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110010011011011010001011100010;
		b = 32'b00111110100011110100001000110010;
		correct = 32'b00110001100001001111101101101111;
		#400 //1.3832251e-08 * 0.2798019 = 3.8702903e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001011011110111111001111000111;
		b = 32'b01010010011100010011101000100010;
		correct = 32'b10011110011011010110100110110101;
		#400 //-4.852424e-32 * 259015600000.0 = -1.2568535e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001110010110101010100111101111;
		b = 32'b01111000001010010001100001100011;
		correct = 32'b11000111000100000110111100000011;
		#400 //-2.6952395e-30 * 1.3718637e+34 = -36975.01
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000101001101110001001110101110;
		b = 32'b10101000100000101100000100001001;
		correct = 32'b00101110001110110000010000010101;
		#400 //-2929.23 * -1.4516615e-14 = 4.2522503e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110010110110110001101010110110;
		b = 32'b01000101111010000001000111111010;
		correct = 32'b01111001010001101001111110011000;
		#400 //8.679617e+30 * 7426.247 = 6.4456983e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101011110111110001101010111110;
		b = 32'b10111110000101100101001110000110;
		correct = 32'b01101010100000110000001001110110;
		#400 //-5.394335e+26 * -0.14680299 = 7.919045e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010010001111111010110011010000;
		b = 32'b01010010010001000101101101011101;
		correct = 32'b01100101000100110000010010110111;
		#400 //205809520000.0 * 210836600000.0 = 4.339218e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110100101001100100010110111000;
		b = 32'b11001000001100110100001110000101;
		correct = 32'b01111101011010001101110100110101;
		#400 //-1.05387615e+32 * -183566.08 = 1.9345592e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001100000010101101111101011101;
		b = 32'b11001111001010011111010100111000;
		correct = 32'b10011011101110000110010011110101;
		#400 //1.0698349e-31 * -2851420200.0 = -3.0505488e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011100101101101001110100100111;
		b = 32'b01000001010101001010011111101111;
		correct = 32'b10011110100101111011000111101111;
		#400 //-1.2084373e-21 * 13.290999 = -1.6061338e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100101110001110101010111001000;
		b = 32'b10100010011001110010001001110111;
		correct = 32'b01001000101100111111100100111110;
		#400 //-1.1766666e+23 * -3.1324583e-18 = 368585.94
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011001100011111100100100000011;
		b = 32'b10110100011100110101001111000011;
		correct = 32'b00001110100010001010101011011010;
		#400 //-1.4867041e-23 * -2.2661611e-07 = 3.3691113e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111100111011101110111000110110;
		b = 32'b01111110001111000001001010100101;
		correct = 32'b11111011101011111000100001010110;
		#400 //-0.029166322 * 6.249792e+37 = -1.8228343e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011111011010001111100110001011;
		b = 32'b00101100111001010011101000010101;
		correct = 32'b10001100110100001001110000010101;
		#400 //-4.9334328e-20 * 6.51502e-12 = -3.2141413e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111010110100101000110101110001;
		b = 32'b00011100001011000001011000011001;
		correct = 32'b01010111100011011000100100110101;
		#400 //5.4662556e+35 * 5.6938587e-22 = 311240880000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011011011011010111000110000001;
		b = 32'b10011000110001000010110000000100;
		correct = 32'b10110100101101011111001110111010;
		#400 //6.683437e+16 * -5.0709257e-24 = -3.3891212e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110111000001111010111001100101;
		b = 32'b00100100100001111110100000110000;
		correct = 32'b00011100000100000001000000001101;
		#400 //8.087231e-06 * 5.894026e-17 = 4.766635e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111110100001001011010011101;
		b = 32'b10100101011011111101101101111101;
		correct = 32'b10101101110000110110111101110011;
		#400 //106797.23 * -2.0804311e-16 = -2.2218427e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011010011110100011000011010010;
		b = 32'b00111001010101111000111100000111;
		correct = 32'b10010100010100101010101011001000;
		#400 //-5.1738225e-23 * 0.0002055728 = -1.0635971e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000011001101010010101100001011;
		b = 32'b10100011001111001000000010011110;
		correct = 32'b10100111000001010110011010100001;
		#400 //181.16814 * -1.0218736e-17 = -1.8513093e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000000000011010101010010110001;
		b = 32'b11101101010111111100101111011111;
		correct = 32'b01101101111101110001101010100111;
		#400 //-2.2082942 * -4.3288514e+27 = 9.559377e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010001001010011011101011111111;
		b = 32'b11001001001101000011100101111010;
		correct = 32'b11011010111011101111101100101110;
		#400 //45561670000.0 * -738199.6 = -3.363361e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000000010110101110101001000111;
		b = 32'b01100000001110001000000001110000;
		correct = 32'b01100001000111011100011000111000;
		#400 //3.4205492 * 5.3178997e+19 = 1.8190137e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001111110011010111100100100000;
		b = 32'b00011000001011000011001110111111;
		correct = 32'b00101000100010100011011011101010;
		#400 //6894534700.0 * 2.2256604e-24 = 1.5344893e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010100110111001010110110111101;
		b = 32'b11100100101111000111101010111001;
		correct = 32'b10111010001000100111100101100001;
		#400 //2.228285e-26 * -2.7814648e+22 = -0.00061978964
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000010111000111010100100101101;
		b = 32'b11000100111001010100010001110001;
		correct = 32'b11001000010010111110001100110011;
		#400 //113.83042 * -1834.1388 = -208780.8
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110001000011110111010001101;
		b = 32'b00010001001000001101111110010010;
		correct = 32'b10000111110010111000010100000111;
		#400 //-2.4129724e-06 * 1.2690667e-28 = -3.0622232e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111011001011011101011011110010;
		b = 32'b00010010101101011000100110110000;
		correct = 32'b10001110011101101000110011110001;
		#400 //-0.0026525822 * 1.14566485e-27 = -3.0389702e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000111011110000101001111001;
		b = 32'b00101101000110010001010100111011;
		correct = 32'b10011110100011101111000100010101;
		#400 //-1.7392515e-09 * 8.701757e-12 = -1.5134544e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010000111110100001101010001000;
		b = 32'b10000000000101000010110100111010;
		correct = 32'b00010000100111011011001000010000;
		#400 //-33568342000.0 * -1.852934e-39 = 6.219993e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010110110110110101110111111;
		b = 32'b10010010011011001100110011101111;
		correct = 32'b00001101110010101111011011111011;
		#400 //-0.0016740485 * -7.472107e-28 = 1.250867e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011100001101110101011000111001;
		b = 32'b11011100001001010100011000010000;
		correct = 32'b01111000111011001011100110000000;
		#400 //-2.064189e+17 * -1.8608162e+17 = 3.8410764e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001110000001110110000100011011;
		b = 32'b01011010010001111001010111110000;
		correct = 32'b01101000110100110001011110001101;
		#400 //567822000.0 * 1.4044595e+16 = 7.97483e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100101100000010001100111011001;
		b = 32'b10111011000100100111001111001000;
		correct = 32'b10100001000100111011011001000010;
		#400 //2.2395448e-16 * -0.0022346843 = -5.0046754e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101000111100011000011011100110;
		b = 32'b01001111001000011001101111111010;
		correct = 32'b01111000100110000111100011111111;
		#400 //9.12463e+24 * 2711353900.0 = 2.47401e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000101101110011010001010001000;
		b = 32'b01100110111101110011101111001001;
		correct = 32'b01101101001100110100011100101011;
		#400 //5940.3164 * 5.8376368e+23 = 3.4677408e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111000011100110111101000011001;
		b = 32'b00001011010110011010100011110001;
		correct = 32'b11000100010011110000001100101101;
		#400 //-1.9753196e+34 * 4.1919777e-32 = -828.0496
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111000001001100111000001111000;
		b = 32'b01110001010101101001000001000100;
		correct = 32'b11101010000010110111111111010000;
		#400 //-3.968223e-05 * 1.0624672e+30 = -4.2161067e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101011111010111101011110100001;
		b = 32'b00100001101001001001111010010100;
		correct = 32'b10001110000101111010100000111011;
		#400 //-1.6757603e-12 * 1.1155048e-18 = -1.8693187e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101100000000110100101010100011;
		b = 32'b00000101000101101101001111110010;
		correct = 32'b10110001100110101011010011011100;
		#400 //-6.34887e+26 * 7.091894e-36 = -4.502551e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010111110001101101010100010010;
		b = 32'b01001100110011111000110100010011;
		correct = 32'b00100101001000010011001111011100;
		#400 //1.2849237e-24 * 108816536.0 = 1.3982095e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010101100100111101010100001101;
		b = 32'b11010111001000100000011110011000;
		correct = 32'b11101101001110110010001001101010;
		#400 //20317907000000.0 * -178153500000000.0 = -3.6197063e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001111011011010000011000110011;
		b = 32'b01000010111110000101011000111111;
		correct = 32'b11010010111001011110110111011100;
		#400 //-3976606500.0 * 124.16845 = -493769060000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010101011100011111001010001100;
		b = 32'b11010100010111010011000010000001;
		correct = 32'b01101010010100010000110000111010;
		#400 //-16626502000000.0 * -3800006100000.0 = 6.318081e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101010111000011111111110001011;
		b = 32'b10011000111101101001000110010100;
		correct = 32'b11000100010110011010110000010100;
		#400 //1.3660754e+26 * -6.3736506e-24 = -870.6887
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111100111011100001110011111011;
		b = 32'b00000111101011111110010111110101;
		correct = 32'b10000101001000111001101110110011;
		#400 //-0.029066553 * 2.646623e-34 = -7.6928206e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010111011000000110111111100010;
		b = 32'b10001011011110111000110100011111;
		correct = 32'b10100011010111001000100101101011;
		#400 //246771140000000.0 * -4.844701e-32 = -1.1955323e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100101000000100011001010010001;
		b = 32'b11000001101010101111101110000111;
		correct = 32'b01100111001011011110101100000001;
		#400 //-3.8427527e+22 * -21.372816 = 8.2130446e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001110110001100011001000111100;
		b = 32'b11101010000010110011100010110000;
		correct = 32'b10111001010101111001001001010100;
		#400 //4.8859142e-30 * -4.2077097e+25 = -0.0002055851
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001100011100011101100011010111;
		b = 32'b01000010101111010100000000001000;
		correct = 32'b00001111101100101100100110010100;
		#400 //1.8631218e-31 * 94.62506 = 1.76298e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110111011101111100011111001010;
		b = 32'b10011100001100001110011111000110;
		correct = 32'b01010100001010110011100110110000;
		#400 //-5.025584e+33 * -5.8533075e-22 = 2941629000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010100010011101101100010001111;
		b = 32'b00110111100001011011001010011000;
		correct = 32'b11001100010110000000110110011111;
		#400 //-3553586000000.0 * 1.5938e-05 = -56637052.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101101000111001110010001100011;
		b = 32'b01000001011001110001111101011001;
		correct = 32'b00101111000011011010010101001100;
		#400 //8.918285e-12 * 14.445153 = 1.28826e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111100100110101110011101101001;
		b = 32'b00111110110001100000101000011010;
		correct = 32'b10111011111011111010101000110000;
		#400 //-0.018909173 * 0.38679582 = -0.007313989
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000110010101000010100001100100;
		b = 32'b10000110111111010101111111011111;
		correct = 32'b10001101110100011111101101011111;
		#400 //13578.098 * -9.530889e-35 = -1.2941135e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100011100110110011101001001011;
		b = 32'b10101100110011001100111001101000;
		correct = 32'b11010000111110000101111100110111;
		#400 //5.7268916e+21 * -5.8209444e-12 = -33335917000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100001010010100111101100110011;
		b = 32'b01001101000010011000110001110011;
		correct = 32'b11101110110110011001011000001001;
		#400 //-2.3344498e+20 * 144230190.0 = -3.3669814e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100100010011011111000010011101;
		b = 32'b00011010000111101000001001110001;
		correct = 32'b00111110111111110000011011100000;
		#400 //1.5195682e+22 * 3.2779004e-23 = 0.49809933
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010100111110100010100000101011;
		b = 32'b01100001110001000011001011010001;
		correct = 32'b01110111001111111011100001101001;
		#400 //8595326000000.0 * 4.5240294e+20 = 3.8885507e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000111011111101000101011001001;
		b = 32'b10111010011010001001010000101100;
		correct = 32'b00000010011001110100000100011010;
		#400 //-1.9149621e-34 * -0.0008872177 = 1.6989883e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010101101111100001001011011011;
		b = 32'b11010010111100010011100111111001;
		correct = 32'b00101001001100110001101011001011;
		#400 //-7.677014e-26 * -518029870000.0 = 3.9769223e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011010000000110110011000001000;
		b = 32'b11011010010110010110111010110011;
		correct = 32'b01110100110111110011010010011101;
		#400 //-9246352000000000.0 * -1.5300446e+16 = 1.4147331e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110001111100100011011011111011;
		b = 32'b00010110000010001001011010101110;
		correct = 32'b01001000100000010011101111000110;
		#400 //2.3987789e+30 * 1.1033539e-25 = 264670.2
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011010110110001111001110110111;
		b = 32'b10001111001011100101100101111011;
		correct = 32'b00101010100100111100000101111011;
		#400 //-3.0533281e+16 * -8.596096e-30 = 2.62467e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011110000010011111100001101111;
		b = 32'b01011100011101000011110101111000;
		correct = 32'b11111011000000111010000111101011;
		#400 //-2.4854546e+18 * 2.7498992e+17 = -6.83475e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101000101100011101111110111111;
		b = 32'b11110011101111011101001010011111;
		correct = 32'b01011101000000111110010010001000;
		#400 //-1.9747982e-14 * -3.0078614e+31 = 5.939919e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111001001000101011011110001101;
		b = 32'b01000001111000000001001000001010;
		correct = 32'b10111011100011100110110000010011;
		#400 //-0.00015517902 * 28.008808 = -0.0043463795
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101101001111101101001111000001;
		b = 32'b01010011001110100000111100000100;
		correct = 32'b11000001000010101011000100001100;
		#400 //-1.0847268e-11 * 799115840000.0 = -8.668224
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110110001100001110001111111101;
		b = 32'b00111001111010110001011011101001;
		correct = 32'b01110000101000100111000100011110;
		#400 //8.969418e+32 * 0.00044839762 = 4.0218658e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001111111000100111111010011011;
		b = 32'b11101000110101010011110100011111;
		correct = 32'b11111001001111001010100101101011;
		#400 //7599896000.0 * -8.0559324e+24 = -6.122425e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100100110010111100111101001111;
		b = 32'b01001010001000101111001000101000;
		correct = 32'b10101111100000011011100111111010;
		#400 //-8.838841e-17 * 2669706.0 = -2.3597108e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001000100001000111110000110011;
		b = 32'b01010101111011000101111100100011;
		correct = 32'b10011110111101001010011101110110;
		#400 //-7.97366e-34 * 32486670000000.0 = -2.5903765e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001111011101000010100100101010;
		b = 32'b11101100010001000101100000110011;
		correct = 32'b00111100001110110100001110100011;
		#400 //-1.2038057e-29 * -9.494639e+26 = 0.0114297
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010100000001101000101100010110;
		b = 32'b01011000110011111101110010110010;
		correct = 32'b11101101010110100111110011101000;
		#400 //-2311436400000.0 * 1828374300000000.0 = -4.226171e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100001000011001010001101000001;
		b = 32'b11010101000100101010101011010011;
		correct = 32'b01110110101000010010010111100111;
		#400 //-1.6214424e+20 * -10078899000000.0 = 1.6342354e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101111111101010010100011100010;
		b = 32'b00001101111011111001010000000110;
		correct = 32'b00111110011001010110111011101100;
		#400 //1.517465e+29 * 1.4765148e-30 = 0.22405595
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111010101111001000000110110100;
		b = 32'b10000101100111100110111001011110;
		correct = 32'b01000000111010010101001010100100;
		#400 //-4.8939125e+35 * -1.4898791e-35 = 7.291338
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111001000001010101001111011001;
		b = 32'b00111101100100011001111000001011;
		correct = 32'b01110111000101111010110110011011;
		#400 //4.3267257e+34 * 0.071102224 = 3.0763983e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101000100110011001100011100111;
		b = 32'b00011100011111010000011101000101;
		correct = 32'b01000101100101111101000001111001;
		#400 //5.802741e+24 * 8.3720074e-22 = 4858.059
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111000000011100111011111011001;
		b = 32'b11000011100111001111001110000100;
		correct = 32'b11111100001011101011000100011011;
		#400 //1.155839e+34 * -313.90247 = -3.628207e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110001100100110101010000001;
		b = 32'b00001001001100110110000011001110;
		correct = 32'b00000111111110100000011111011111;
		#400 //0.1742344 * 2.1591859e-33 = 3.7620445e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111001010100010010111001011010;
		b = 32'b00101110101110000000000001111110;
		correct = 32'b11101000100101100101100110111000;
		#400 //-6.7883135e+34 * 8.367439e-11 = -5.68008e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111110011100001001111011001010;
		b = 32'b01000001101101101001100011101100;
		correct = 32'b11000000101010111010000010100000;
		#400 //-0.23498073 * 22.824669 = -5.3633575
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101000101101100110111001110000;
		b = 32'b00110111100000100000001101000010;
		correct = 32'b00100000101110010100110011001110;
		#400 //2.0253954e-14 * 1.5498725e-05 = 3.1391044e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010110100000101010011011100100;
		b = 32'b11011110001001000001111101100101;
		correct = 32'b00110101001001111000010111100000;
		#400 //-2.1107956e-25 * -2.9565705e+18 = 6.240716e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000010001011010000110000100001;
		b = 32'b11101000110011110111001010000100;
		correct = 32'b00101011100011000011101000110111;
		#400 //-1.2713513e-37 * -7.8371384e+24 = 9.963756e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100000111010001000110000001001;
		b = 32'b10100111011011101001101101001001;
		correct = 32'b11001000110110001011111100111111;
		#400 //1.3405423e+20 * -3.3113315e-15 = -443897.97
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000010110000111100001100100000;
		b = 32'b01111011111010101011011101111110;
		correct = 32'b00111111001100110111110010101100;
		#400 //2.876467e-37 * 2.4374383e+36 = 0.7011211
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011011101101101100100111111000;
		b = 32'b10000101110101101101011101100011;
		correct = 32'b10100010000110010110011010100000;
		#400 //1.02901026e+17 * -2.0203584e-35 = -2.0789696e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110011011001111011011011011010;
		b = 32'b11011100110100001011110110101101;
		correct = 32'b01010000101111001111000001000000;
		#400 //-5.395018e-08 * -4.7004277e+17 = 25358893000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101101000000010111001011101110;
		b = 32'b01011101001110001010010001010011;
		correct = 32'b01001010101110101011101101100101;
		#400 //7.3583206e-12 * 8.3155315e+17 = 6118834.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011110011010101100011000000001;
		b = 32'b01101000010010000110100100101111;
		correct = 32'b01000111001101111100101100100111;
		#400 //1.2428803e-20 * 3.7856544e+24 = 47051.152
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111000111011001101101010011000;
		b = 32'b11010011011010111001101001011100;
		correct = 32'b01001100110110011111101101111010;
		#400 //-0.00011294073 * -1011907040000.0 = 114285520.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000000111010000001100101000011;
		b = 32'b11011000101000111010011011110110;
		correct = 32'b10011010000101000101111101110101;
		#400 //2.1314897e-38 * -1439499900000000.0 = -3.0682792e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111111110001001010110100111111;
		b = 32'b11001111000100001111001001101101;
		correct = 32'b11001111010111101011011101100110;
		#400 //1.536537 * -2431806700.0 = -3736561200.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100101101000000101101000010010;
		b = 32'b00011111110101110100000110001110;
		correct = 32'b01000110000001101101010010110101;
		#400 //9.465502e+22 * 9.116449e-20 = 8629.177
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001000010000001010111001111011;
		b = 32'b01101100111101000010110001010000;
		correct = 32'b00110101101101111100011110100111;
		#400 //5.7983e-34 * 2.3614973e+27 = 1.3692669e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000001010100011010001001001000;
		b = 32'b01000110101111101110111010110101;
		correct = 32'b00001000100111000101100111101011;
		#400 //3.8503668e-38 * 24439.354 = 9.410048e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000010101101110010000100111011;
		b = 32'b00110001110011100100011111110110;
		correct = 32'b10110101000100111001000000111000;
		#400 //-91.5649 * 6.00357e-09 = -5.4971633e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100010000101111100001011001011;
		b = 32'b01001011100100100111110001111111;
		correct = 32'b01101110001011011010110111001011;
		#400 //6.998737e+20 * 19200254.0 = 1.3437752e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111000101000001000101100111101;
		b = 32'b00000101011111111100001110110010;
		correct = 32'b00111110101000000110010101101011;
		#400 //2.6049737e+34 * 1.2025986e-35 = 0.31327376
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011000010110001110001110110010;
		b = 32'b10111001101001111100111111000000;
		correct = 32'b01010010100011100010110010001100;
		#400 //-953889800000000.0 * -0.00032007508 = 305316360000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011101001100110010011111100000;
		b = 32'b11100000110000000100010010101011;
		correct = 32'b00111110100001101000110111110110;
		#400 //-2.3711068e-21 * -1.1083509e+20 = 0.26280183
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000001101101110000101111110100;
		b = 32'b00011100011101101111010001010111;
		correct = 32'b00011110101100001001010000110010;
		#400 //22.880836 * 8.1710374e-22 = 1.8696017e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110100101000010110010010111111;
		b = 32'b11010010110010001111000101111011;
		correct = 32'b11000111111111010101110111100101;
		#400 //3.006189e-07 * -431522400000.0 = -129723.79
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001100111110001101101001101110;
		b = 32'b10110110000100001110101011111000;
		correct = 32'b11000011100011001101111101000111;
		#400 //130470770.0 * -2.1594442e-06 = -281.74435
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100001101001011000001100111000;
		b = 32'b11011001111100000000010110100001;
		correct = 32'b00111100000110110010111010101000;
		#400 //-1.1215568e-18 * -8445023000000000.0 = 0.009471573
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011001000000001000010101000110;
		b = 32'b01000010010100100001010110001010;
		correct = 32'b01011011110100101111000001000111;
		#400 //2260958300000000.0 * 52.521034 = 1.18747866e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111111011110001001000110000;
		b = 32'b01000100000111110001010010101101;
		correct = 32'b01001100100101001000111110011011;
		#400 //122404.375 * 636.32306 = 77888730.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111000111001010110111001010111;
		b = 32'b11111100001011100111111100010010;
		correct = 32'b01110101100111000110001011100001;
		#400 //-0.00010940123 * -3.6241478e+36 = 3.9648624e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000001100100000101101101100100;
		b = 32'b01001000001011010100001000011111;
		correct = 32'b00001010010000110110011000010111;
		#400 //5.3028385e-38 * 177416.48 = 9.4081094e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000101101100101010100001100111;
		b = 32'b01000001001101011011111001010000;
		correct = 32'b11000111011111011010101111000011;
		#400 //-5717.0503 * 11.358963 = -64939.76
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101100001111111100101100101101;
		b = 32'b01010101001011110110101001110110;
		correct = 32'b11000010000000110110101110100110;
		#400 //-2.7255518e-12 * 12054486000000.0 = -32.855125
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101101101011001010111000100101;
		b = 32'b10110100000111111001010010010001;
		correct = 32'b00100010010101110100100010111111;
		#400 //-1.9631472e-11 * -1.4862077e-07 = 2.9176445e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010110000101011000111101111111;
		b = 32'b11111011111011011101010101011100;
		correct = 32'b01010010100010101111001001111111;
		#400 //-1.2081404e-25 * -2.4698036e+36 = 298386950000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010100001000001001000001011100;
		b = 32'b01011010101011001100100110101111;
		correct = 32'b10101111010110001011111011111010;
		#400 //-8.1064055e-27 * 2.4317725e+16 = -1.9712934e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100011101000111111110000110110;
		b = 32'b00100111101011011111111100011001;
		correct = 32'b11001011110111101110100110110001;
		#400 //-6.049986e+21 * 4.8293723e-15 = -29217634.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111011101110111001101010011111;
		b = 32'b11000011010110000001011011010010;
		correct = 32'b00111111100111100101101100101111;
		#400 //-0.0057252194 * -216.08914 = 1.2371577
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101111100000111100011011111110;
		b = 32'b01101100011101011110100000100011;
		correct = 32'b11011100011111010010100111011111;
		#400 //-2.3970154e-10 * 1.18913224e+27 = -2.8503683e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011011000001100010001100011111;
		b = 32'b00101111001100111000110000100011;
		correct = 32'b00001010101111000010011111111000;
		#400 //1.1095568e-22 * 1.6329742e-10 = 1.8118776e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101111111001101001110000110011;
		b = 32'b01001000100011101010000001010100;
		correct = 32'b01111001000000000111101100010010;
		#400 //1.4274077e+29 * 292098.62 = 4.1694385e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010100001000110111111101111101;
		b = 32'b10000011100110101100110001001011;
		correct = 32'b10011000010001011011101001010101;
		#400 //2808874300000.0 * -9.09821e-37 = -2.5555727e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101010000100100001000000111101;
		b = 32'b10111111101110100110111101111101;
		correct = 32'b11101010010101001011111011010001;
		#400 //4.4144963e+25 * -1.4565274 = -6.4298345e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011101010000101001011100101110;
		b = 32'b00101110101001100010000110111000;
		correct = 32'b01001100011111001000111101010010;
		#400 //8.763579e+17 * 7.554796e-11 = 66207050.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110010111000110101101001100010;
		b = 32'b00111111111000101101111100001101;
		correct = 32'b10110011010010010111101111100010;
		#400 //-2.646738e-08 * 1.772432 = -4.691163e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010001110110111101001010101000;
		b = 32'b11101011110110011001100110100110;
		correct = 32'b11111110001110101101100110000000;
		#400 //118016510000.0 * -5.2612497e+26 = -6.2091433e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101010000000101111101110000000;
		b = 32'b10010110010110100111100010001101;
		correct = 32'b10000000110111111000111110110010;
		#400 //1.1633576e-13 * -1.7647939e-25 = -2.0530864e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111011011100111001011001010101;
		b = 32'b01000100111001010100010111101001;
		correct = 32'b11000000110110100010011111111111;
		#400 //-0.0037168462 * 1834.1847 = -6.8173823
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100101101110110100101100010101;
		b = 32'b10011011001010010011101011011000;
		correct = 32'b10000001011101111001111100111100;
		#400 //3.2490207e-16 * -1.3998366e-22 = -4.548098e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001111101001011011000000000010;
		b = 32'b11000000101000101001000010010100;
		correct = 32'b00010000110100100110110111101000;
		#400 //-1.6338052e-29 * -5.0801487 = 8.299973e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100111001111001000111110000110;
		b = 32'b01000110000010010000010101010011;
		correct = 32'b11101101110010011101100101110101;
		#400 //-8.9045244e+23 * 8769.331 = -7.808672e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000101111100010111010110111111;
		b = 32'b11110111111000000101000011011010;
		correct = 32'b10111110010100111001001101001010;
		#400 //2.2706784e-35 * -9.099331e+33 = -0.20661655
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111001111101010100111101110001;
		b = 32'b00001100000011010110101111111010;
		correct = 32'b11000110100001111000010000111001;
		#400 //-1.592155e+35 * 1.0894738e-31 = -17346.111
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011110110101001100101011011110;
		b = 32'b01101010101000010110100010110110;
		correct = 32'b11001010000001100010101010011111;
		#400 //-2.2530277e-20 * 9.756577e+25 = -2198183.8
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000100010010010001010110010101;
		b = 32'b11010000100111110101101011111110;
		correct = 32'b10010101011110100101011111000001;
		#400 //2.3637346e-36 * -21388325000.0 = -5.0556324e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011011010000101011110000000;
		b = 32'b00001110011100110101100110011111;
		correct = 32'b10011010010111001101110001100101;
		#400 //-15226752.0 * 2.9995213e-30 = -4.5672967e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001101000011000011011011000101;
		b = 32'b01000110010111011000010101111100;
		correct = 32'b01010011111100101010100011001001;
		#400 //147024980.0 * 14177.371 = 2084427700000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101111110010011000100100000100;
		b = 32'b01010100011000110000111011100110;
		correct = 32'b01000100101100101100000000111001;
		#400 //3.6659042e-10 * 3900830000000.0 = 1430.007
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111101111110100010111001000100;
		b = 32'b00110010010110011001010001000110;
		correct = 32'b00110000110101001010001000011111;
		#400 //0.12215856 * 1.2664776e-08 = 1.5471108e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110011110000010110000101100110;
		b = 32'b11111101011111001000000101100010;
		correct = 32'b11110001101111101011110110011101;
		#400 //9.0049795e-08 * -2.0977328e+37 = -1.8890042e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100010010110001010101011100001;
		b = 32'b00111011111100000110010111001101;
		correct = 32'b00011110110010110111011001011100;
		#400 //2.9363921e-18 * 0.0073363543 = 2.1542413e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011111100110010011100010000010;
		b = 32'b01011100000011001000101111100111;
		correct = 32'b11111100001010000011110101000110;
		#400 //-2.2081435e+19 * 1.5824128e+17 = -3.4941946e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100000000100000111000001011000;
		b = 32'b11010000111000010100100111010111;
		correct = 32'b01110001011111100011100011001101;
		#400 //-4.163166e+19 * -30237702000.0 = 1.2588458e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011001000001110100101000010111;
		b = 32'b01101001101100111110000011110010;
		correct = 32'b11000011001111100001111101011110;
		#400 //-6.994299e-24 * 2.71825e+25 = -190.12253
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111100001001110111100101110001;
		b = 32'b01001001101000111001100011011100;
		correct = 32'b11000110010101100000110010100110;
		#400 //-0.010221825 * 1340187.5 = -13699.162
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101011010010011101111001100101;
		b = 32'b00111000111010001001110000011001;
		correct = 32'b01100100101101110110110010100011;
		#400 //2.4404432e+26 * 0.000110916975 = 2.7068658e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101101111001011100010110011001;
		b = 32'b11011101110011100010101110010101;
		correct = 32'b01001100001110010000110000011111;
		#400 //-2.6122037e-11 * -1.8570165e+18 = 48509052.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101000111010000010011100010100;
		b = 32'b11000101100011000101001111011100;
		correct = 32'b11101110111111101000001011010110;
		#400 //8.770479e+24 * -4490.4824 = -3.9383682e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001000110101110111100110010000;
		b = 32'b00111111010010010100100001001010;
		correct = 32'b11001000101010010110101101001011;
		#400 //-441292.5 * 0.7862593 = -346970.34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110011100101111101001100000101;
		b = 32'b11111011101100011101010101011110;
		correct = 32'b01101111110100101110111011100010;
		#400 //-7.06987e-08 * -1.8467283e+36 = 1.3056129e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101000100010001011001011111010;
		b = 32'b11000010111011111011010100011001;
		correct = 32'b10101011111111111111111110010111;
		#400 //1.5176652e-14 * -119.85371 = -1.818978e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010100100010110010100100001010;
		b = 32'b01001011001110000101010011011011;
		correct = 32'b00100000010010000110011100111111;
		#400 //1.40516e-26 * 12080347.0 = 1.697482e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011000100011000001000101111010;
		b = 32'b11010100111111011011100000110000;
		correct = 32'b01101110000010101101001000001100;
		#400 //-1232053500000000.0 * -8717735000000.0 = 1.0740716e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001001001110011001000000101000;
		b = 32'b00111001000000111101011111000101;
		correct = 32'b10000010101111110010001001010111;
		#400 //-2.2336347e-33 * 0.00012573514 = -2.8084638e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111100110011010101101111101001;
		b = 32'b10010111010001100010110001011110;
		correct = 32'b00010100100111101111100010101101;
		#400 //-0.02506824 * -6.403325e-25 = 1.6052008e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111100010010000111000010110101;
		b = 32'b00011011110100110011010011101100;
		correct = 32'b11011000101001010101111001010101;
		#400 //-4.1629814e+36 * 3.4941222e-22 = -1454596600000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101100111100010000011111110100;
		b = 32'b10101010011000101111100010010110;
		correct = 32'b01010111110101011011001100010010;
		#400 //-2.3311094e+27 * -2.0159078e-13 = 469930160000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100000111001000001101100000000;
		b = 32'b11001000011001000111100110111010;
		correct = 32'b10101001110010111001010010000010;
		#400 //3.864257e-19 * -233958.9 = -9.040773e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010100110110010001100100010000;
		b = 32'b01110110111001111011001001110111;
		correct = 32'b11001100010001000111110011110110;
		#400 //-2.1921286e-26 * 2.349688e+33 = -51508184.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111111011011111110011100011101;
		b = 32'b00101000100010100101100100011001;
		correct = 32'b00101000100000011010011000010100;
		#400 //0.93712026 * 1.5359718e-14 = 1.4393902e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000000100010110011001110001001;
		b = 32'b01100111001101010010101111100010;
		correct = 32'b01101000010001010000011010011001;
		#400 //4.350041 * 8.555578e+23 = 3.7217116e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000101101011000010001011001101;
		b = 32'b11100000111100010101100010000101;
		correct = 32'b00100111001000100100100001001000;
		#400 //-1.6187586e-35 * -1.3912637e+20 = 2.25212e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011100101101000011010001010110;
		b = 32'b00011110001110110010111000101101;
		correct = 32'b10111011100000111100001010111100;
		#400 //-4.0578432e+17 * 9.9092465e-21 = -0.004021017
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011111011101100101011111100000;
		b = 32'b10100110011110001000110111011011;
		correct = 32'b11000110011011110010110110100010;
		#400 //1.7750903e+19 * -8.6234534e-16 = -15307.408
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101111000010010000000111101010;
		b = 32'b10100011111000110101001001010001;
		correct = 32'b01010011011100110101000110000001;
		#400 //-4.240176e+28 * -2.4646252e-17 = 1045044460000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101111101010011001100101101000;
		b = 32'b01010111010011100010101101101110;
		correct = 32'b01000111100010001001011000110111;
		#400 //3.0849923e-10 * 226685920000000.0 = 69932.43
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100111010100010111111011011000;
		b = 32'b10101100100101111000000000100000;
		correct = 32'b00010100011101111111010101010110;
		#400 //-2.9073339e-15 * -4.305903e-12 = 1.2518697e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010001000100111111110101000110;
		b = 32'b11010011110000111110110001010001;
		correct = 32'b11100101011000101000010100010001;
		#400 //39725590000.0 * -1682966700000.0 = -6.685684e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100010100010010011010110011000;
		b = 32'b10001111101010001011001001110001;
		correct = 32'b10110010101101001101010110011111;
		#400 //1.2655329e+21 * -1.6634812e-29 = -2.1051902e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000011001010101001001100100101;
		b = 32'b00010000110110111011110101011011;
		correct = 32'b10010100100100100110101000001100;
		#400 //-170.57478 * 8.667202e-29 = -1.478406e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010010000111110010011111001000;
		b = 32'b01011101001001011001100111110011;
		correct = 32'b11101111110011011110100010110100;
		#400 //-170891800000.0 * 7.4580224e+17 = -1.274515e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000010111101001001110111111110;
		b = 32'b11000110101001101110100000000110;
		correct = 32'b11001010000111110111110000101000;
		#400 //122.30858 * -21364.012 = -2613002.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011111101000101101010111101011;
		b = 32'b00100010111001100010111001110011;
		correct = 32'b01000011000100100110100110111101;
		#400 //2.3467086e+19 * 6.2390805e-18 = 146.41304
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101000111011011011110001011110;
		b = 32'b00011000100000011111110000010101;
		correct = 32'b11000001111100010110110000001001;
		#400 //-8.981405e+24 * 3.3600256e-24 = -30.177752
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101110111111110000110000011011;
		b = 32'b01010000111010111000010000110110;
		correct = 32'b11000000011010101010001111010101;
		#400 //-1.1598208e-10 * 31610483000.0 = -3.6662495
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100010000110011111110110111000;
		b = 32'b00101001110000111110011100101111;
		correct = 32'b11001100011010111010111010100111;
		#400 //-7.1015855e+20 * 8.6998436e-14 = -61782684.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110111010001001000100100000001;
		b = 32'b11010011001110000000111100110111;
		correct = 32'b11001011000011010100111000100111;
		#400 //1.1714409e-05 * -790529250000.0 = -9260583.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001110011010100000010101001111;
		b = 32'b10110111100011011100000001011100;
		correct = 32'b10000110100000011001010011000101;
		#400 //2.8845283e-30 * -1.6898084e-05 = -4.8743004e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111111100101001010011100111101;
		b = 32'b00011110100010011000000110011110;
		correct = 32'b10011110100111111011000110000111;
		#400 //-1.1613537 * 1.4559048e-20 = -1.6908203e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010111110110101001100001010101;
		b = 32'b10111001101000101001110101111101;
		correct = 32'b10010010000010101101101011100000;
		#400 //1.4126374e-24 * -0.00031016386 = -4.3814906e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000011110010101111011111100;
		b = 32'b01011011000101111001111011101011;
		correct = 32'b11001100000100111011000111010100;
		#400 //-9.0720653e-10 * 4.2677454e+16 = -38717264.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101110101110100000110101100100;
		b = 32'b10110101010101010011101100000011;
		correct = 32'b10100100100110101111100000000111;
		#400 //8.4606794e-11 * -7.9434557e-07 = -6.720703e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001111000001110111000110000001;
		b = 32'b11110110101101111111010100101111;
		correct = 32'b11000110010000101010011110110111;
		#400 //6.677874e-30 * -1.8655532e+33 = -12457.929
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000101010001010101110001110100;
		b = 32'b01100010011000011000011111001011;
		correct = 32'b01101000001011011101111011110010;
		#400 //3157.7783 * 1.0400756e+21 = 3.284328e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011001110000100000010011011100;
		b = 32'b01000101001001111111110001001100;
		correct = 32'b01011111011111101010000011000100;
		#400 //6826436000000000.0 * 2687.7686 = 1.834788e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010110001111111011001001001;
		b = 32'b11101100101111011000101101000011;
		correct = 32'b01101000000101000000110110011011;
		#400 //-0.0015255894 * -1.833157e+27 = 2.796645e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110011101111011100100000100100;
		b = 32'b10001111111111001011010000010111;
		correct = 32'b11000100001110110101011010000101;
		#400 //3.0072126e+31 * -2.4918487e-29 = -749.35187
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111101000100000001100101111110;
		b = 32'b11001111000111001111010000100110;
		correct = 32'b11001100101100001011000111101101;
		#400 //0.03518056 * -2633246200.0 = -92639080.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110001110010011101011100011001;
		b = 32'b01110101111100011000011011100011;
		correct = 32'b11101000001111100110110111011000;
		#400 //-5.8743237e-09 * 6.1234344e+32 = -3.5971036e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111000101100110001010001000101;
		b = 32'b01101101111001100101001100100111;
		correct = 32'b01100111001000010001111001100001;
		#400 //8.5391606e-05 * 8.9102597e+27 = 7.608614e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111001011100101000011000010010;
		b = 32'b00010100011000110101100010011011;
		correct = 32'b01001110010101110110000011010011;
		#400 //7.8703444e+34 * 1.14780456e-26 = 903361700.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001100111010100011001001000000;
		b = 32'b11010100111000111011100110010011;
		correct = 32'b00100010010100000101010001010100;
		#400 //-3.6083652e-31 * -7824568000000.0 = 2.82339e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001101111100110100111101010111;
		b = 32'b10010110010010111111110101101101;
		correct = 32'b10100100110000011110000011000111;
		#400 //510257900.0 * -1.6478176e-25 = -8.4081195e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011101011101010110001010000000;
		b = 32'b01111111111111011100010010001010;
		correct = 32'b01111111111111011100010010001010;
		#400 //3.2476403e-21 * nan = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101001111011010100101111001000;
		b = 32'b11000011000101111110000011100010;
		correct = 32'b10101101100011001100100000100111;
		#400 //1.053806e-13 * -151.87845 = -1.6005043e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101111011010100100110011010101;
		b = 32'b00101100010010011001001010011011;
		correct = 32'b11011100001110000111110010000001;
		#400 //-7.2512377e+28 * 2.86452e-12 = -2.0771316e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001011000011010001101011111110;
		b = 32'b11001011111001010100000101110010;
		correct = 32'b00010111011111001011101001110000;
		#400 //-2.717592e-32 * -30048996.0 = 8.166091e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000110100011000111010000010100;
		b = 32'b00010000111100000111100001011100;
		correct = 32'b00011000000000111110111011011100;
		#400 //17978.04 * 9.484875e-29 = 1.7051946e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100111000000001011001000111010;
		b = 32'b11100001001111010111110111111111;
		correct = 32'b01001000101111101000010111011000;
		#400 //-1.7860185e-15 * -2.184696e+20 = 390190.75
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100010101000001110100011110100;
		b = 32'b11111011111000011100110001111110;
		correct = 32'b11011111000011011110110101000111;
		#400 //4.3614736e-18 * -2.3448288e+36 = -1.0226908e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001101001001010100010100110100;
		b = 32'b11010100001110000110001110010000;
		correct = 32'b01100001111011100001010000001000;
		#400 //-173298500.0 * -3167777500000.0 = 5.4897106e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000101011100111101001010111000;
		b = 32'b11001100100010000000001010000000;
		correct = 32'b10010010100000011000101001010011;
		#400 //1.1464508e-35 * -71308290.0 = -8.175144e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010101000011101000000010010011;
		b = 32'b00111001000111100011010011000110;
		correct = 32'b11001110101100000010000101110110;
		#400 //-9792680000000.0 * 0.00015087714 = -1477491500.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101001101000111111010001011110;
		b = 32'b10111001111101111100001000110000;
		correct = 32'b01100100000111101010110100100101;
		#400 //-2.4776113e+25 * -0.00047256192 = 1.1708248e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000101101000111100110101111001;
		b = 32'b01100011111100101010101101000101;
		correct = 32'b10101010000110110100010111010011;
		#400 //-1.5403925e-35 * 8.9529067e+21 = -1.379099e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110101001101111100011110010010;
		b = 32'b01011111101011100100110000010110;
		correct = 32'b11010101011110100100000010001001;
		#400 //-6.8463225e-07 * 2.5118875e+19 = -17197193000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001100001011011000110101111011;
		b = 32'b11111001101101010001001100111100;
		correct = 32'b01000110011101011000010000100100;
		#400 //-1.337001e-31 * -1.1752448e+35 = 15713.035
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101110110111011111001001110110;
		b = 32'b11100000101010001001010001100011;
		correct = 32'b11010000000100100010011111000011;
		#400 //1.0092986e-10 * -9.717954e+19 = -9808317000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010100000011111010101000000011;
		b = 32'b10100000100010010000110110010110;
		correct = 32'b10110101000110011101001100110111;
		#400 //2468130600000.0 * -2.3217693e-19 = -5.73043e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110101101110111000111111000;
		b = 32'b10100101010101011110011011110000;
		correct = 32'b00011100100110010100011101010000;
		#400 //-5.4670927e-06 * -1.855305e-16 = 1.0143125e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000101100101001001011100001110;
		b = 32'b11000101100101111010010010001000;
		correct = 32'b01001011101100000000100100110010;
		#400 //-4754.882 * -4852.5664 = 23073380.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110010001011101110101111011111;
		b = 32'b01011000101001011111111111000010;
		correct = 32'b01001011011000101101100110010000;
		#400 //1.0181764e-08 * 1460143100000000.0 = 14866832.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111011011101010111010110111110;
		b = 32'b01010011011111001100100110011010;
		correct = 32'b11001111011100100110000100110100;
		#400 //-0.0037454213 * 1085714100000.0 = -4066456600.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111001111011001011100000101001;
		b = 32'b01011100011000111000111110110001;
		correct = 32'b01010110110100100110110000101011;
		#400 //0.00045150638 * 2.5621124e+17 = 115681010000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011010000001010100110011111011;
		b = 32'b11010100110000011101110111010111;
		correct = 32'b11101111010010011110010100011001;
		#400 //9380203000000000.0 * -6661204300000.0 = -6.248345e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001000001001110110001111001010;
		b = 32'b10111001011011011101011111101011;
		correct = 32'b01000010000110111000010010010000;
		#400 //-171407.16 * -0.00022682517 = 38.879456
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111111011110110000110110110010;
		b = 32'b10111101000110111000101011011101;
		correct = 32'b11111101000110001000100101111001;
		#400 //3.3370734e+38 * -0.037974227 = -1.2672278e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011100000110000011100111100110;
		b = 32'b00011101110111100001100101100110;
		correct = 32'b00111010100001000001000101010000;
		#400 //1.7139143e+17 * 5.8789172e-21 = 0.001007596
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111011111111101110100100111111;
		b = 32'b01010001000001000001011010001110;
		correct = 32'b11001101100000111000011010111010;
		#400 //-0.00777927 * 35457130000.0 = -275830600.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110011110111010001001100100101;
		b = 32'b01011101001000100111011111000010;
		correct = 32'b01010001100011000100110110001001;
		#400 //1.0294597e-07 * 7.3168994e+17 = 75324530000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111110101110111011011010010001;
		b = 32'b10100001011100011001001000111101;
		correct = 32'b00100000101100010010001000011001;
		#400 //-0.36662725 * -8.184752e-19 = 3.000753e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110011111111101000111111110;
		b = 32'b01001100001000101100110100000010;
		correct = 32'b01001011001000101010111111000000;
		#400 //0.2498245 * 42677256.0 = 10661824.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001001011110110001110010111101;
		b = 32'b01100101100101011111000001100110;
		correct = 32'b10101111100100110001001110001001;
		#400 //-3.0226539e-33 * 8.85084e+22 = -2.6753025e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110111101011110100100000110101;
		b = 32'b10110001001000010000001110100100;
		correct = 32'b10101001010111000111110111001111;
		#400 //2.089525e-05 * -2.3430653e-09 = -4.8958935e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100001010001110100110110100000;
		b = 32'b10100111100101000110101110011000;
		correct = 32'b00001001011001110001100101001001;
		#400 //-6.752656e-19 * -4.1194905e-15 = 2.7817503e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110001000011001010011110001010;
		b = 32'b00101010100001100011111010000001;
		correct = 32'b11011100000100111000010000010011;
		#400 //-6.964871e+29 * 2.3846552e-13 = -1.6608815e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001111100110100110100001111100;
		b = 32'b00011111111110011000010101001101;
		correct = 32'b00110000000101101000000000000111;
		#400 //5181077500.0 * 1.0567613e-19 = 5.475162e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111111001101011010011000111010;
		b = 32'b10001101000010010110010001010101;
		correct = 32'b01001100110000101111101001001101;
		#400 //-2.4145336e+38 * -4.2337155e-31 = 102224490.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111000001100011111100101000110;
		b = 32'b00010100100001110111001101001000;
		correct = 32'b10001101001111000101010100110010;
		#400 //-4.2432242e-05 * 1.3676987e-26 = -5.8034523e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111101001110101110101011000101;
		b = 32'b00111110000010111100111111100001;
		correct = 32'b10111011110011000010101010000010;
		#400 //-0.04563405 * 0.13653518 = -0.0062306533
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100010001010001001110000101001;
		b = 32'b11101110101110010100110010001111;
		correct = 32'b11010001011101000001011010001100;
		#400 //2.2850916e-18 * -2.867364e+28 = -65521893000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111001110000000101001110110001;
		b = 32'b00111010111011000101111101001011;
		correct = 32'b11110101001100011001010010111111;
		#400 //-1.2482731e+35 * 0.0018033771 = -2.2511071e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000111010010110001110011110;
		b = 32'b10011111010110001101000111001010;
		correct = 32'b00010000110001011010101101010000;
		#400 //-1.6981294e-09 * -4.5913313e-20 = 7.796675e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001100011000101010011101101101;
		b = 32'b00110111011111010110001000101100;
		correct = 32'b11000100011000000101011001100010;
		#400 //-59415988.0 * 1.5102833e-05 = -897.34973
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011011011101000110110000110100;
		b = 32'b01010000001011111101100000100000;
		correct = 32'b00101100001001111110010001010001;
		#400 //2.0218169e-22 * 11800707000.0 = 2.3858868e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110101000010100001000111100001;
		b = 32'b00100100100100101101100101001011;
		correct = 32'b11011010000111100110011011001000;
		#400 //-1.7502431e+32 * 6.3685515e-17 = -1.1146514e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101000000011100110011100101011;
		b = 32'b11001100101110010100010000000010;
		correct = 32'b00110101010011100001110011000101;
		#400 //-7.9049545e-15 * -97132560.0 = 7.6782845e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110001010011111101000010111100;
		b = 32'b01000111110101010001001100110001;
		correct = 32'b00111001101011001111100001000001;
		#400 //3.0241116e-09 * 109094.38 = 0.0003299136
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100110101100001101010110110000;
		b = 32'b11010010011000010110001001001001;
		correct = 32'b01111001100110111010111110110100;
		#400 //-4.1753917e+23 * -242004150000.0 = 1.0104621e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000001111111101101110011000101;
		b = 32'b10100100010110100000111110001001;
		correct = 32'b00100110110110010001011101110111;
		#400 //-31.857798 * -4.7284374e-17 = 1.506376e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110100001111100000101101011100;
		b = 32'b00001101011000001101000010110011;
		correct = 32'b01000010001001101110010011011111;
		#400 //6.0227466e+31 * 6.927654e-31 = 41.723507
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010110000110100110010101010000;
		b = 32'b10001110100110101111001100111011;
		correct = 32'b00100101001110101110011101001000;
		#400 //-42439980000000.0 * -3.8198153e-30 = 1.621129e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011010010010000101100001110100;
		b = 32'b10110010011001011000111101001011;
		correct = 32'b01001101001100111010011101000100;
		#400 //-1.4098063e+16 * -1.3362135e-08 = 188380220.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101111111111100010010111001101;
		b = 32'b00010010111111001011011001010110;
		correct = 32'b10000011011110101110001000111010;
		#400 //-4.622919e-10 * 1.5948385e-27 = -7.3728092e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100001001111100010111111100101;
		b = 32'b00100011101011000000011010101001;
		correct = 32'b10000101011111111001101001000001;
		#400 //-6.443789e-19 * 1.8651098e-17 = -1.2018374e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010000000001010100011011011100;
		b = 32'b01100101111000101001110000100101;
		correct = 32'b01110110011010111111001110110001;
		#400 //8944054000.0 * 1.337669e+23 = 1.1964184e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111101101110000010100110010110;
		b = 32'b10010010010001011100101101010100;
		correct = 32'b00010000100011100100101001000110;
		#400 //-0.08992307 * -6.241286e-28 = 5.612356e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110001010100010001110010000101;
		b = 32'b11001101010010010111101110111001;
		correct = 32'b11111111001001001001010001110100;
		#400 //1.0354695e+30 * -211270540.0 = -2.187642e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001111000000000000110000001110;
		b = 32'b00111110110100010001111111110000;
		correct = 32'b00001110010100010011001110100010;
		#400 //6.313209e-30 * 0.4084468 = 2.57861e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110111001011010000111110000010;
		b = 32'b00000011101100000011011010111101;
		correct = 32'b10111011011011100011111101010101;
		#400 //-3.5100855e+33 * 1.0356918e-36 = -0.0036353667
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111010100110010001010100101;
		b = 32'b01011000100100011000110110100101;
		correct = 32'b11010000011100000001011011100011;
		#400 //-1.2584646e-05 * 1280300400000000.0 = -16112127000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101100010111111101001100101101;
		b = 32'b10010100000000100001011000001110;
		correct = 32'b10000000111000110111100100001010;
		#400 //3.1807432e-12 * -6.567672e-27 = -2.0890078e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110111010101010000000000101;
		b = 32'b00101111101011111100010101101101;
		correct = 32'b00101111001000010001100001010100;
		#400 //0.4582521 * 3.1972594e-10 = 1.4651508e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110010100111010011100111100101;
		b = 32'b10101011001111100000010101011111;
		correct = 32'b11011110011010010110100010001001;
		#400 //6.2283695e+30 * -6.7509014e-13 = -4.2047109e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111011100101100101001100110111;
		b = 32'b10001111000100100110110001011010;
		correct = 32'b01001011001010111111011000101011;
		#400 //-1.5610647e+36 * -7.2192235e-30 = 11269675.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101111111100010101100111111000;
		b = 32'b00100111111001110100100100110010;
		correct = 32'b10011000010110100000110100110001;
		#400 //-4.390157e-10 * 6.419474e-15 = -2.81825e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100000110011100101011100010010;
		b = 32'b00101110001011000001111010111100;
		correct = 32'b00001111100010101011101101000110;
		#400 //3.4955376e-19 * 3.913557e-11 = 1.3679986e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111110111100000011110110100111;
		b = 32'b10011010001111110110101011110010;
		correct = 32'b00011001101100111010001001011100;
		#400 //-0.46922037 * -3.9584264e-23 = 1.8573743e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110101100001101101111101010011;
		b = 32'b11100010101100000000011000110101;
		correct = 32'b11011000101110010111100110011100;
		#400 //1.0048774e-06 * -1.6235371e+21 = -1631455700000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101010000100110110111110001011;
		b = 32'b10000001100110011100111010110011;
		correct = 32'b10101100001100010010100101101010;
		#400 //4.455971e+25 * -5.649992e-38 = -2.5176202e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010100001101010101010101010010;
		b = 32'b00011000001100101110111100100011;
		correct = 32'b10101100111111010111110101101101;
		#400 //-3115282000000.0 * 2.3126694e-24 = -7.2046175e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000001110101000001111110001010;
		b = 32'b01011001000100111111101111100011;
		correct = 32'b11011011011101010011110110100111;
		#400 //-26.5154 * 2603361000000000.0 = -6.9029157e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111010100011110010010110111001;
		b = 32'b10001010101011100101100110110101;
		correct = 32'b11000101110000101111101110011010;
		#400 //3.7163178e+35 * -1.6789335e-32 = -6239.45
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101111111010111110000000101101;
		b = 32'b01001001111111001110010100011100;
		correct = 32'b00111010011010010000001111000110;
		#400 //4.2905537e-10 * 2071715.5 = 0.0008888807
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011111000011101011010110001100;
		b = 32'b01011101010000100000110000100000;
		correct = 32'b10111100110110000101100010101101;
		#400 //-3.0219842e-20 * 8.739116e+17 = -0.026409471
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011011111001010010011010101101;
		b = 32'b01101111011101101100010011001100;
		correct = 32'b01001011110111001110001101010010;
		#400 //3.7909866e-22 * 7.6371225e+28 = 28952228.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000100011011101101001011010010;
		b = 32'b11100100100001001110111101100111;
		correct = 32'b00101001011110000000100000010110;
		#400 //-2.807357e-36 * -1.9617768e+22 = 5.5074075e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111001010000010111010000001110;
		b = 32'b00111110110010001101010001000110;
		correct = 32'b10111000100101111100001100010100;
		#400 //-0.00018449148 * 0.39224452 = -7.236577e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011001111001110101101110111110;
		b = 32'b10010100100100111101001111100000;
		correct = 32'b00101111000001011001100100101001;
		#400 //-8140199000000000.0 * -1.4926777e-26 = 1.2150693e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110110110110111011010010010010;
		b = 32'b00100101101100111011010111100011;
		correct = 32'b11011101000110100011101101011100;
		#400 //-2.228077e+33 * 3.1174801e-16 = -6.945986e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101000100111110010010011101000;
		b = 32'b10111011011101100001011010000110;
		correct = 32'b10100100100110001111101101110111;
		#400 //1.7668552e-14 * -0.0037550046 = -6.634549e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110100000000101000100000000110;
		b = 32'b11011111101001001001011101111111;
		correct = 32'b11010100001001111101100011000110;
		#400 //1.2156679e-07 * -2.3720176e+19 = -2883585600000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101101001100100111001101010100;
		b = 32'b11100111011010101010101000101110;
		correct = 32'b11010101001000111001010000001011;
		#400 //1.01437365e-11 * -1.108173e+24 = -11241015000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110101100000000110111001000001;
		b = 32'b10100011110110110110111001010111;
		correct = 32'b01011001110111000010101101011001;
		#400 //-3.2561046e+32 * -2.3790758e-17 = 7746519500000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110010110110010110101000000111;
		b = 32'b10001100011100101001111000110111;
		correct = 32'b10111111110011100000110010011001;
		#400 //8.6126626e+30 * -1.8690613e-31 = -1.6097594
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101101001000110100101100001001;
		b = 32'b11010101101010001010000010000000;
		correct = 32'b11000011010101110001111100111101;
		#400 //9.282138e-12 * -23175912000000.0 = -215.12202
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111100001110001001110110001110;
		b = 32'b11100101101010011100111001010001;
		correct = 32'b11100010011101001110100110011000;
		#400 //0.011268033 * -1.00235725e+23 = -1.12945944e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000111010010100001110001010010;
		b = 32'b01100010101011110111101010001100;
		correct = 32'b10101010100010101000101000011100;
		#400 //-1.5205114e-34 * 1.6185053e+21 = -2.4609557e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100101010100000000101111111000;
		b = 32'b01000100110110011011011001111010;
		correct = 32'b10101010101100001110111001110001;
		#400 //-1.8045179e-16 * 1741.7024 = -3.1429332e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001011110010011110101100111111;
		b = 32'b01110100101100011000100011100000;
		correct = 32'b01000001000011000000011110011100;
		#400 //7.777634e-32 * 1.1252596e+32 = 8.751858
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101001101001001110001001000110;
		b = 32'b10100001110101011111111110001000;
		correct = 32'b01001100000010011101010011011001;
		#400 //-2.4916548e+25 * -1.450108e-18 = 36131684.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101000000111110001010101010000;
		b = 32'b10000111101101111001100100011001;
		correct = 32'b00110000011001000010111010111111;
		#400 //-3.0049977e+24 * -2.7624762e-34 = 8.3012347e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000000000101110010111000101110;
		b = 32'b11000001100111110111010100000110;
		correct = 32'b00000001011001110000010001110100;
		#400 //-2.128783e-39 * -19.93214 = 4.2431194e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100000011011110110110100000;
		b = 32'b10111010011001010111000011000000;
		correct = 32'b10111110111111100110100000100101;
		#400 //567.7129 * -0.0008752458 = -0.4968883
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110100100010111001111100001;
		b = 32'b11010011111111100000100100000110;
		correct = 32'b11010011000100000101011000011010;
		#400 //0.2840872 * -2182146200000.0 = -619919840000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000000000001000000001100111010;
		b = 32'b11100100011110001010111110100000;
		correct = 32'b01100101000000000011110110110001;
		#400 //-2.062697 * -1.8349791e+22 = 3.7850057e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001011101010101001100101111000;
		b = 32'b11001101110110011111110111000110;
		correct = 32'b10011010000100010100010100110100;
		#400 //6.571253e-32 * -457160900.0 = -3.00412e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110101100001010001100011001010;
		b = 32'b01010111101110101110000100110001;
		correct = 32'b01001101110000100101001000101110;
		#400 //9.916487e-07 * 410952700000000.0 = 407520700.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010111110001001100011111100001;
		b = 32'b11000110011000010100010100100101;
		correct = 32'b01011110101011010010100011010011;
		#400 //-432725500000000.0 * -14417.286 = 6.2387274e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011011000010010110000100000100;
		b = 32'b00111000111100111011011000100111;
		correct = 32'b10010100100000101100100011010111;
		#400 //-1.1363722e-22 * 0.000116210715 = -1.3205863e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101000011010010010111011101010;
		b = 32'b00110000001001100000101011010100;
		correct = 32'b10011001000101110011111001001001;
		#400 //-1.2944271e-14 * 6.0405836e-10 = -7.8190954e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001010110010010011010000101010;
		b = 32'b11100000000110111101010100001110;
		correct = 32'b11101011011101001111010000010010;
		#400 //6593045.0 * -4.4915587e+19 = -2.9613049e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100110101001101011110001110001;
		b = 32'b00000000001011010010001110110101;
		correct = 32'b00100110111010110011001100001100;
		#400 //3.936945e+23 * 4.145407e-39 = 1.6320237e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011011010001011100110010010111;
		b = 32'b00111100010100101101011110110010;
		correct = 32'b00011000001000101110100001111100;
		#400 //1.6361565e-22 * 0.012868809 = 2.1055384e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101101010001000110101110010011;
		b = 32'b10010011001000010110000101111011;
		correct = 32'b00000000111101111010010011100101;
		#400 //-1.1165196e-11 * -2.0369119e-27 = 2.274252e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001101100111011011010001111010;
		b = 32'b10000101110011110101000000001101;
		correct = 32'b00010011111111110110110001111110;
		#400 //-330731330.0 * -1.9495592e-35 = 6.447803e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110101100001111010010111001100;
		b = 32'b10110011001011011101111101011010;
		correct = 32'b10101001001110000100001011001000;
		#400 //1.0106537e-06 * -4.048284e-08 = -4.091413e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011011101010100100001110001110;
		b = 32'b11000101100100001100011011111110;
		correct = 32'b10100001110000001001010010110010;
		#400 //2.8167797e-22 * -4632.874 = -1.3049785e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100110000110100011100011100101;
		b = 32'b11001110010010011000110101000010;
		correct = 32'b11110100111100101101011110001010;
		#400 //1.8207349e+23 * -845369500.0 = -1.5391937e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100010010110000010010001111101;
		b = 32'b01000110110101010001100010101001;
		correct = 32'b10101001101100111110101100101110;
		#400 //-2.9292775e-18 * 27276.33 = -7.989994e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001010010000111011101001010000;
		b = 32'b10010111100101111010111001010100;
		correct = 32'b10100010011001111111000001011100;
		#400 //3206804.0 * -9.802153e-25 = -3.1433583e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100010001000010010010101000000;
		b = 32'b00100010010111001000000100011100;
		correct = 32'b00000101000010101100110101001000;
		#400 //2.1839289e-18 * 2.988391e-18 = 6.526433e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011100101101000000000111011111;
		b = 32'b01110100110101001111001100010110;
		correct = 32'b11010010000101011011110001111010;
		#400 //-1.1911884e-21 * 1.3497282e+32 = -160778060000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000011010100010000001110110001;
		b = 32'b00001110001100000001011000100001;
		correct = 32'b00010010000011111100010010011011;
		#400 //209.01442 * 2.170433e-30 = 4.536518e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101000100101110101111111101000;
		b = 32'b11011111001100010101010000101100;
		correct = 32'b11001000010100011011011000101010;
		#400 //1.680596e-14 * -1.2777886e+19 = -214744.66
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101000001110101011010000000001;
		b = 32'b10110110001100100010001110101111;
		correct = 32'b10011111000000011110101100101111;
		#400 //1.0364106e-14 * -2.6544838e-06 = -2.7511352e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000111101010010000110001010101;
		b = 32'b01011101100100011101100110010110;
		correct = 32'b11100101110000001001111101010101;
		#400 //-86552.664 * 1.3136995e+18 = -1.1370419e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111110110001001000010100110011;
		b = 32'b10011000000001010100010000101100;
		correct = 32'b11010111010011001001101100010001;
		#400 //1.3061015e+38 * -1.7224265e-24 = -224966380000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001111111101111010101100010110;
		b = 32'b10100010011001011011010100100101;
		correct = 32'b00110010110111100011101101001010;
		#400 //-8310369300.0 * -3.1131184e-18 = 2.5871163e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111111111011111000000101011110;
		b = 32'b11011001000001101000000110010111;
		correct = 32'b11111111111011111000000101011110;
		#400 //nan * -2366258300000000.0 = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101111101011110110011001000111;
		b = 32'b11000000111010000100010101000001;
		correct = 32'b10110001000111110010010000100011;
		#400 //3.1904987e-10 * -7.258454 = -2.3158087e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100000001000010001101101000110;
		b = 32'b10101000011100100100000100100100;
		correct = 32'b01001001000110000111010011000111;
		#400 //-4.6435798e+19 * -1.3447824e-14 = 624460.44
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100111110100001010011000110001;
		b = 32'b10100011010110010000111111110100;
		correct = 32'b10001011101100001110100111100000;
		#400 //5.7911782e-15 * -1.1766972e-17 = -6.814463e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101111100110011101010101101010;
		b = 32'b00011100001100011011011010011111;
		correct = 32'b11001100010101011001010010010111;
		#400 //-9.521842e+28 * 5.880042e-22 = -55988828.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001100111011000000100010011011;
		b = 32'b11110000101010100100000010000000;
		correct = 32'b10111110000111001111100100101111;
		#400 //3.6366737e-31 * -4.2152342e+29 = -0.15329431
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001111110111011010000111011000;
		b = 32'b10010001001111101111110110101110;
		correct = 32'b10100001101001010101100110111110;
		#400 //7436742700.0 * -1.5066528e-28 = -1.1204589e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011011111100001101110110111101;
		b = 32'b01010101110001010000010000011010;
		correct = 32'b10110010001110010101111001111110;
		#400 //-3.9847964e-22 * 27077676000000.0 = -1.0789902e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000110010000001010011000111010;
		b = 32'b01001010111111101101011111111111;
		correct = 32'b11010001101111111100011101111001;
		#400 //-12329.557 * 8350719.5 = -102960670000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110001010101100001101110011110;
		b = 32'b10101101100101010110111000001011;
		correct = 32'b00011111011110011111010000111000;
		#400 //-3.1156797e-09 * -1.6988208e-11 = 5.2929814e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101110110100010110011001101010;
		b = 32'b00111001101101001010001010010000;
		correct = 32'b11101001000100111100000011111011;
		#400 //-3.240309e+28 * 0.00034453394 = -1.1163964e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111011010011000100100000111110;
		b = 32'b10100001100111111001011111011001;
		correct = 32'b00011101011111101011010000010101;
		#400 //-0.003117099 * -1.0814453e-18 = 3.370972e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001000110011000000000111110011;
		b = 32'b01101010111110111111001000100011;
		correct = 32'b11110100010010001100011011011111;
		#400 //-417807.6 * 1.5229192e+26 = -6.362872e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111101010100100111001100000;
		b = 32'b00101010111111001011011010110111;
		correct = 32'b00110011001010000001111010110100;
		#400 //87196.75 * 4.4890976e-13 = 3.9143472e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000011010001010000101010000001;
		b = 32'b11101001001101001010101101101100;
		correct = 32'b00101101000010110000111101010100;
		#400 //-5.7905155e-37 * -1.365101e+25 = 7.904639e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010001010011101100110101111111;
		b = 32'b11100110010000001011101100110001;
		correct = 32'b10111000000110111011000101010111;
		#400 //1.6313858e-28 * -2.2753686e+23 = -3.712004e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010110001110011011011011111011;
		b = 32'b00011000111100111010101111010011;
		correct = 32'b00101111101100001100010101010111;
		#400 //51048887000000.0 * 6.2987526e-24 = 3.2154432e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100100110011101001110100101100;
		b = 32'b11101100101100110111000010111101;
		correct = 32'b01010010000100001101001011100011;
		#400 //-8.960452e-17 * -1.7354409e+27 = 155503350000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101010000001001011110110110100;
		b = 32'b01101010001001101011011001100100;
		correct = 32'b11010100101011001110001100101011;
		#400 //-1.1789772e-13 * 5.038575e+25 = -5940365000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101101111101111100010110000011;
		b = 32'b10101010111000011101010110000111;
		correct = 32'b11011001010110101001001101000010;
		#400 //9.585197e+27 * -4.0116193e-13 = -3845216000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000011000101010001001111111000;
		b = 32'b00001110001000000101001010000111;
		correct = 32'b10010001101110101011100100010100;
		#400 //-149.078 * 1.9761258e-30 = -2.945969e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010111101010010001100000100011;
		b = 32'b11011000010011010101100010110110;
		correct = 32'b00110000100001111010001011101101;
		#400 //-1.0927462e-24 * -903123600000000.0 = 9.868849e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110100010011010000111111000001;
		b = 32'b00101111011000000101111010010111;
		correct = 32'b10100100001100111011100110001110;
		#400 //-1.9097844e-07 * 2.0406286e-10 = -3.897161e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000000000100010010001110101101;
		b = 32'b11101110011100100110000000011001;
		correct = 32'b01101111000010010110101000110101;
		#400 //-2.2678025 * -1.8752887e+28 = 4.2527843e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101100010000110010011101100001;
		b = 32'b00100101001110010100101111100000;
		correct = 32'b11010010000011010100000101001100;
		#400 //-9.43706e+26 * 1.60719e-16 = -151671470000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100101111111101101010001110010;
		b = 32'b01000100101100000011101010100000;
		correct = 32'b10101011001011110110110001101010;
		#400 //-4.4205935e-16 * 1409.832 = -6.2322944e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010110001110101100001000100111;
		b = 32'b00000011111011000001000001000000;
		correct = 32'b10011010101011000011011011010111;
		#400 //-51335760000000.0 * 1.3874564e-36 = -7.122613e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111100001001101101011011000000;
		b = 32'b10111000000110010001000111011111;
		correct = 32'b10110100110001111000001111111101;
		#400 //0.010183036 * -3.6494686e-05 = -3.7162673e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010000100011001100010110001010;
		b = 32'b01001100000001100001110101010110;
		correct = 32'b00011101000100110111111100010000;
		#400 //5.552462e-29 * 35157336.0 = 1.9520978e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011100111011010100000001011010;
		b = 32'b01011100100010111000101111001001;
		correct = 32'b01111010000000010101001101111101;
		#400 //5.342426e+17 * 3.1422974e+17 = 1.678749e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000010100000101001101011010010;
		b = 32'b10001000000101011111101111011101;
		correct = 32'b00001011000110010000100100110110;
		#400 //-65.30238 * -4.513412e-34 = 2.9473658e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011111100111100110101010101101;
		b = 32'b00001000000111100110101110111001;
		correct = 32'b00101000010001000001000100000000;
		#400 //2.2830253e+19 * 4.7673023e-34 = 1.0883872e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100111011110100111100101011100;
		b = 32'b01111101001101001011111001101110;
		correct = 32'b01100101001100001101011110100110;
		#400 //3.4760259e-15 * 1.5015613e+37 = 5.2194657e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110111010111100001000011001010;
		b = 32'b11010010010001000100101001110100;
		correct = 32'b11001010001010100100010101110000;
		#400 //1.323614e-05 * -210765680000.0 = -2789724.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001110001100111011111011110100;
		b = 32'b11111000110010110101010011001001;
		correct = 32'b01000111100011101100001111110011;
		#400 //-2.2155394e-30 * -3.2992372e+34 = 73095.9
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010101101100111001011011111111;
		b = 32'b11101110001100000110001011000110;
		correct = 32'b11000100011101110111101000110100;
		#400 //7.2535754e-26 * -1.3647193e+28 = -989.9094
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101110001101000011011100010110;
		b = 32'b00111010010000110111000100111110;
		correct = 32'b10101001000010011001010110101110;
		#400 //-4.0976188e-11 * 0.0007455534 = -3.0549937e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000000100111000000011100111110;
		b = 32'b10101000100000100101100101011000;
		correct = 32'b10101001100111101110010001000011;
		#400 //4.875884 * -1.4471646e-14 = -7.0562066e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111100111010100101111101011110;
		b = 32'b00001110010111011010001100011111;
		correct = 32'b00001011110010101110100110101011;
		#400 //0.028609928 * 2.7318893e-30 = 7.8159154e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101111101101111111001111001111;
		b = 32'b10100000110100111111101011010011;
		correct = 32'b01010001000110000101001000101111;
		#400 //-1.1386101e+29 * -3.5910772e-19 = 40888365000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111100001001010101100011000100;
		b = 32'b11110001001110111010000110101011;
		correct = 32'b01101101111100100110000010000101;
		#400 //-0.010091964 * -9.291063e+29 = 9.376507e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110101100001110111100010111;
		b = 32'b10011011011011100000010000101001;
		correct = 32'b10011010101001001000000100100111;
		#400 //0.3455741 * -1.9688243e-22 = -6.803747e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000111011110111110110001111111;
		b = 32'b11100111100100001111100100011100;
		correct = 32'b00101111100011101010101000101100;
		#400 //-1.8952641e-34 * -1.369232e+24 = 2.5950564e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100001101101100011100101100000;
		b = 32'b00101110111000000011011110100000;
		correct = 32'b10010001000111111001100111001100;
		#400 //-1.2347987e-18 * 1.01962216e-10 = -1.2590281e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011000000110001010110010100100;
		b = 32'b01011000000011101100100111100010;
		correct = 32'b01110000101010100101000001010011;
		#400 //671469000000000.0 * 627990900000000.0 = 4.2167646e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111100110010110100001111000001;
		b = 32'b10101001011110111000100001110001;
		correct = 32'b00100110110001111011011111000100;
		#400 //-0.024812581 * -5.585154e-14 = 1.3858209e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010010000001101011001101010;
		b = 32'b11110111101111000010000001000101;
		correct = 32'b01110010100011011011010111000101;
		#400 //-0.0007356169 * -7.6312993e+33 = 5.613713e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100100010110111000000011111111;
		b = 32'b11110110111110011100000111000001;
		correct = 32'b11011011110101100010011010011010;
		#400 //4.759732e-17 * -2.5328354e+33 = -1.2055618e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001000010001101101011110010001;
		b = 32'b01001000110001010010011011111100;
		correct = 32'b00010001100110010010001000101010;
		#400 //5.9836855e-34 * 403767.88 = 2.41602e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100000110101001010001000010000;
		b = 32'b10111000011001000001000111101010;
		correct = 32'b01011001101111010110111100110111;
		#400 //-1.2257461e+20 * -5.437612e-05 = 6665131600000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110100011111001001010000001100;
		b = 32'b10100100010101001100101110001011;
		correct = 32'b01011001010100011111001101101100;
		#400 //-8.004526e+31 * -4.614258e-17 = 3693494700000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001010110100001100110011110000;
		b = 32'b10100000111000011101100011010110;
		correct = 32'b00101100001110000011010011111010;
		#400 //-6841976.0 * -3.8259973e-19 = 2.617738e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111110101011111000110100010111;
		b = 32'b00111101000111011101001110001011;
		correct = 32'b10111100010110000111010100101111;
		#400 //-0.3428733 * 0.03853182 = -0.0132115325
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011000001000001101000011011010;
		b = 32'b11000011111100011001000010100010;
		correct = 32'b01011100100101111011111101111000;
		#400 //-707275500000000.0 * -483.12994 = 3.4170595e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001111110001001101100001100110;
		b = 32'b00000110100100100111100101100101;
		correct = 32'b00010110111000010100000110000100;
		#400 //6605032400.0 * 5.509747e-35 = 3.6392057e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000110110111000011101101011001;
		b = 32'b01101011000010110101010001000110;
		correct = 32'b11110010011011111011100101110010;
		#400 //-28189.674 * 1.6843866e+26 = -4.7482308e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011010111101110110111111101110;
		b = 32'b11110000110011000100100100000111;
		correct = 32'b11001100010001010111001111000111;
		#400 //1.0233764e-22 * -5.057858e+29 = -51760924.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010110111000100000100001011111;
		b = 32'b10011110110000111010011101011000;
		correct = 32'b00110110001011001100000000100010;
		#400 //-124262790000000.0 * -2.071564e-20 = 2.5741833e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011011101010011011110101110010;
		b = 32'b10110100010100110101010111101100;
		correct = 32'b11010000100011000010000000011101;
		#400 //9.555514e+16 * -1.9682165e-07 = -18807319000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110011111000100001000100100011;
		b = 32'b01100100100101010111111100100111;
		correct = 32'b11011001000001000000010001000010;
		#400 //-1.0527062e-07 * 2.2061817e+22 = -2322461200000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001011000111110100000111000111;
		b = 32'b11000100111011101111111000011010;
		correct = 32'b11010000100101001010110100111010;
		#400 //10437063.0 * -1911.9407 = -19955044000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100110001100010000011000110011;
		b = 32'b00011001000101001000100101000001;
		correct = 32'b00111111110011010110110011111101;
		#400 //2.089933e+23 * 7.679139e-24 = 1.6048886
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100110110010010001101110000101;
		b = 32'b01101100001100010101001100000001;
		correct = 32'b01010011100010110100110100111100;
		#400 //1.3954636e-15 * 8.574874e+26 = 1196592500000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101110001010000101101001101010;
		b = 32'b11010000010101001101110011110100;
		correct = 32'b01111111000010111111110000101110;
		#400 //-1.3025696e+28 * -14285001000.0 = 1.8607208e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001110000110100001110110110000;
		b = 32'b10001101011011111000011100111001;
		correct = 32'b10011100000100000011001100011111;
		#400 //646409200.0 * -7.381033e-31 = -4.7711676e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100111011010111001111010010010;
		b = 32'b10010000001110010010101100000101;
		correct = 32'b10111000001010100110110100110000;
		#400 //1.1126812e+24 * -3.6517958e-29 = -4.0632847e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000000001100110110000110100011;
		b = 32'b11010101101100101100011100111100;
		correct = 32'b11010110011110101000101011111101;
		#400 //2.8028343 * -24571097000000.0 = -68868714000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111001111101101010000000100100;
		b = 32'b01011010010010011101010001101101;
		correct = 32'b01010100110000100111000001100010;
		#400 //0.0004704009 * 1.4202509e+16 = 6680873000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111000000110000010010000111001;
		b = 32'b10100100001010111011111110011100;
		correct = 32'b00011100110011000010010000100100;
		#400 //-3.627336e-05 * -3.7242014e-17 = 1.350893e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110001011111001000101011100110;
		b = 32'b00111111100001101011001101000101;
		correct = 32'b00110001100001001110000110001110;
		#400 //3.674978e-09 * 1.0523459 = 3.867348e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001101111110101001110011110010;
		b = 32'b01110101000000000000001011010001;
		correct = 32'b11000011011110101010001001110110;
		#400 //-1.5445223e-30 * 1.6227322e+32 = -250.63461
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000110011000110010101001010011;
		b = 32'b01000110110011000110111000000101;
		correct = 32'b11001101101101010110011101011011;
		#400 //-14538.581 * 26167.01 = -380431200.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000111101011111100111100001000;
		b = 32'b00111000110001001100110010110000;
		correct = 32'b10000001000001110010011100010100;
		#400 //-2.6452755e-34 * 9.384134e-05 = -2.482362e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110001111110101000010010000;
		b = 32'b00101100010011010110010110110001;
		correct = 32'b10100011000110010111111110000010;
		#400 //-2.8508111e-06 * 2.9188702e-12 = -8.3211474e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100100011010111000100111010111;
		b = 32'b10110110000100111100111000011001;
		correct = 32'b00011011000001111111110111000110;
		#400 //-5.1074257e-17 * -2.2024672e-06 = 1.1248937e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011000100100010110111010010110;
		b = 32'b00010100111001001001101001010100;
		correct = 32'b10101110000000011101111000101010;
		#400 //-1279233200000000.0 * 2.3082988e-26 = -2.9528525e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110001010110011011101010111110;
		b = 32'b10001111010110111011111001011110;
		correct = 32'b00000001001110101110010010101001;
		#400 //-3.1683807e-09 * -1.0834197e-29 = 3.432686e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100100011100000111100110110110;
		b = 32'b00100111110010000011001000101100;
		correct = 32'b10001100101111000000111000110111;
		#400 //-5.2144797e-17 * 5.5565548e-15 = -2.8974542e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110001110010110010011111010111;
		b = 32'b01010110011100110001100000001001;
		correct = 32'b01001000110000001110100111100100;
		#400 //5.912607e-09 * 66821140000000.0 = 395087.12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100111110101011100000001011101;
		b = 32'b11001101011111000111010111001101;
		correct = 32'b01110101110100101100101110111000;
		#400 //-2.0188251e+24 * -264723660.0 = 5.344308e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110101110001100111111001001101;
		b = 32'b11010011101010010111000001011000;
		correct = 32'b11001010000000110110000001111100;
		#400 //1.4788908e-06 * -1455468600000.0 = -2152479.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110101000110101011100100000101;
		b = 32'b11010010011001111101010101010011;
		correct = 32'b11001000000011000001110111100010;
		#400 //5.763871e-07 * -248929100000.0 = -143479.53
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000010010001110011101101010001;
		b = 32'b01001101001011111001100101100011;
		correct = 32'b01010000000010001010100011101100;
		#400 //49.807926 * 184129070.0 = 9171087000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000111000100111100001111111101;
		b = 32'b00010110010100100100010001101010;
		correct = 32'b10011101111100101011110010000110;
		#400 //-37827.99 * 1.6985253e-25 = -6.4251795e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100111001110011110000111101100;
		b = 32'b00101111101001000100110000000000;
		correct = 32'b01010111011011101001011111010101;
		#400 //8.778053e+23 * 2.9885427e-10 = 262335880000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010011001110110000100011100000;
		b = 32'b00011100101110001000110001010100;
		correct = 32'b00110000100001101101010011100111;
		#400 //803307800000.0 * 1.2212373e-21 = 9.810294e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000010001011010010110101101011;
		b = 32'b01001000110001001110000001000011;
		correct = 32'b00001011100001010010111001111011;
		#400 //1.2723067e-37 * 403202.1 = 5.129967e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011000011111010101101011101010;
		b = 32'b11100010111000111111111101110001;
		correct = 32'b01111011111000011010010001101011;
		#400 //-1114267660000000.0 * -2.1029087e+21 = 2.3432032e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110111110001010000111010000100;
		b = 32'b11001100011001101001101101111100;
		correct = 32'b11000100101100011000001010111010;
		#400 //2.349099e-05 * -60452336.0 = -1420.0852
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110100000011100110110010000001;
		b = 32'b10110011000000101110000000010100;
		correct = 32'b11100111100100011001111110000111;
		#400 //4.513592e+31 * -3.047178e-08 = -1.3753718e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100100111111000011111011001111;
		b = 32'b10111100100101010111110000011101;
		correct = 32'b11100010000100110100101011011001;
		#400 //3.7224843e+22 * -0.018247658 = -6.792662e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010101111100100111101110001111;
		b = 32'b00110000111111110100001110001000;
		correct = 32'b11000111011100011100100100001011;
		#400 //-33326562000000.0 * 1.8572885e-09 = -61897.043
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001100001100011011010110001110;
		b = 32'b00011110110110010110111000001111;
		correct = 32'b00101011100101101110111101001100;
		#400 //46585400.0 * 2.3021288e-20 = 1.0724559e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010001000001111010011111110010;
		b = 32'b01101100111010100100101010111001;
		correct = 32'b01111110011110000100111000111000;
		#400 //36414890000.0 * 2.2659321e+27 = 8.251367e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010011111100000011000001101001;
		b = 32'b01101001111001111001011011111111;
		correct = 32'b00111110010110010100100101011010;
		#400 //6.0632254e-27 * 3.4996865e+25 = 0.21219388
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111110101010110000010101001;
		b = 32'b00111111010101100010001000110010;
		correct = 32'b10110111101100100111101101001110;
		#400 //-2.543659e-05 * 0.8364593 = -2.1276672e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111001111011011111010110111100;
		b = 32'b00111000111000110111110010011100;
		correct = 32'b11110011010100110111010010111010;
		#400 //-1.5444481e+35 * 0.00010847414 = -1.6753267e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100000110101111110100101000101;
		b = 32'b11010111100111110000001000011010;
		correct = 32'b01111001000001100001101110101000;
		#400 //-1.2446434e+20 * -349662750000000.0 = 4.3520545e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001101011100001011110101010110;
		b = 32'b01100110010001000101001011111110;
		correct = 32'b11110100001110001001111100000001;
		#400 //-252433760.0 * 2.317787e+23 = -5.8508765e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010100010100110000011101100111;
		b = 32'b11011100111010110101000011101011;
		correct = 32'b11110001110000011111101010000000;
		#400 //3625449200000.0 * -5.2988472e+17 = -1.9210702e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111111011000000111101101000011;
		b = 32'b11111011001100001010110101110110;
		correct = 32'b11111011000110101110110011011001;
		#400 //0.8768808 * -9.1736245e+35 = -8.0441756e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010001001110100010101010001100;
		b = 32'b11010011101110100110110001111011;
		correct = 32'b01100101100001111001000111001101;
		#400 //-49973610000.0 * -1601367800000.0 = 8.002613e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100101110111111111110001110011;
		b = 32'b10101111100001100101101000000000;
		correct = 32'b10010101111010110001100111000110;
		#400 //3.88554e-16 * -2.4438407e-10 = -9.495641e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100110011100001001000010000101;
		b = 32'b00001100100001010100110101011111;
		correct = 32'b10110011011110101000011110010100;
		#400 //-2.8400847e+23 * 2.053846e-31 = -5.833097e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100000111010010110000111100110;
		b = 32'b01110010000100101111110011011010;
		correct = 32'b01010011100001100000000001011000;
		#400 //3.953652e-19 * 2.9113914e+30 = 1151062800000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000000001001100010111101010000;
		b = 32'b00010011011101010100100101111000;
		correct = 32'b00010100000111110011101011111001;
		#400 //2.5966377 * 3.095957e-27 = 8.039079e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010100001001001010010110110010;
		b = 32'b01011100011010100011001111011001;
		correct = 32'b00110001000101101010000011001101;
		#400 //8.312562e-27 * 2.636886e+17 = 2.1919278e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100001100100111000010010101000;
		b = 32'b10101011101101011101001111010101;
		correct = 32'b01001101110100011000110110111000;
		#400 //-3.401538e+20 * -1.2919619e-12 = 439465730.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000010101001010011001001001010;
		b = 32'b10110010001010111101100110001111;
		correct = 32'b00110101010111011100100111110111;
		#400 //-82.59822 * -1.0002977e-08 = 8.2622813e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011010101010001001000011000101;
		b = 32'b01011111110010001111000001100100;
		correct = 32'b01111011000001000100111101100011;
		#400 //2.3723486e+16 * 2.8958366e+19 = 6.869933e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110011010010110100000110110;
		b = 32'b11111111011010101110100000100101;
		correct = 32'b01110110010101100010110011101010;
		#400 //-3.4780364e-06 * -3.1224471e+38 = 1.0859985e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011001110101001011000100001100;
		b = 32'b10000100010111001111110111101011;
		correct = 32'b00011110101101111001101100011101;
		#400 //-7483420000000000.0 * -2.597747e-36 = 1.9440032e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001000011011101111110011110100;
		b = 32'b11001111001000100110110001010010;
		correct = 32'b10011000000101111010000100110010;
		#400 //7.1917865e-34 * -2725008000.0 = -1.9597675e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001110011110011001001011110111;
		b = 32'b11001101010010001111010101100110;
		correct = 32'b11011100010000111110101000001110;
		#400 //1046789570.0 * -210720350.0 = -2.2057987e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000010100100000010010101000011;
		b = 32'b10011000111111000010000101100010;
		correct = 32'b10011100000011011111011101111010;
		#400 //72.07278 * -6.517418e-24 = -4.697284e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000110001101000011010101101001;
		b = 32'b11110010011110011000111011001000;
		correct = 32'b00111001001011111010110001110110;
		#400 //-3.3893477e-35 * -4.9430003e+30 = 0.00016753547
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010101101001101110111000000111;
		b = 32'b10001011011101101100010110101010;
		correct = 32'b00100001101000001110100110011111;
		#400 //-22942656000000.0 * -4.7526583e-32 = 1.0903861e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001010011000011111000111111100;
		b = 32'b11110011101110011111100100011000;
		correct = 32'b00111110101001000010001110111001;
		#400 //-1.0878868e-32 * -2.9468602e+31 = 0.32058504
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000000000100001001000010001000;
		b = 32'b01000101010100110101001110101110;
		correct = 32'b00000100110110101100100010100011;
		#400 //1.521216e-39 * 3381.23 = 5.143581e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100001010110110111111000010101;
		b = 32'b01110010011110001000000011110111;
		correct = 32'b01010100010101010001000010110111;
		#400 //7.4366954e-19 * 4.9221242e+30 = 3660433900000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010111111111001111011001111;
		b = 32'b01001001001001111001101000101111;
		correct = 32'b11000100101001110101101010001101;
		#400 //-0.0019502285 * 686498.94 = -1338.8297
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111101110010101011011110000111;
		b = 32'b10001101001110010000001011000011;
		correct = 32'b11001011100100101000000011010000;
		#400 //3.3682123e+37 * -5.701085e-31 = -19202464.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101001011100100010110100101010;
		b = 32'b11000110100001000001010001011111;
		correct = 32'b11110000011110011110010100011110;
		#400 //1.8298333e+25 * -16906.186 = -3.0935501e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000001110001000010011010111010;
		b = 32'b00110010111001100101011111101010;
		correct = 32'b00110101001100000111111000101000;
		#400 //24.51891 * 2.6815503e-08 = 6.574869e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101110001001101110110111110100;
		b = 32'b11010101011111111010100000010101;
		correct = 32'b01000100001001101011010010100000;
		#400 //-3.7955375e-11 * -17568586000000.0 = 666.82227
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011011110010111001001110010111;
		b = 32'b10110000101101001110101010111110;
		correct = 32'b00001101000011111101111001110010;
		#400 //-3.367891e-22 * -1.3163441e-09 = 4.4333036e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010000001001101000010110100000;
		b = 32'b10111111001100011111100110100011;
		correct = 32'b01001111111001111000100110001011;
		#400 //-11175100000.0 * -0.6952154 = 7769102000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101100101011111100001101010110;
		b = 32'b00001111010010001011000101101000;
		correct = 32'b10111100100010011100101001101001;
		#400 //-1.6998757e+27 * 9.8949285e-30 = -0.01682015
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111110011010011011001111010;
		b = 32'b00011010011101011101100100010001;
		correct = 32'b00100010110001010001001100100100;
		#400 //105068.95 * 5.0840157e-23 = 5.3417223e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110100101010111011000001100;
		b = 32'b10000100011110000100100100010110;
		correct = 32'b10000011100100001111010100000111;
		#400 //0.29191625 * -2.918582e-36 = -8.519815e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010001000101111010110011110111;
		b = 32'b10000011110101110101001010111101;
		correct = 32'b10010101011111110010011010010010;
		#400 //40715120000.0 * -1.265556e-36 = -5.1527267e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001100010010110000011100100100;
		b = 32'b01010011111111111111111010101101;
		correct = 32'b11100000110010110000011000010111;
		#400 //-53222544.0 * 2198978800000.0 = -1.1703525e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011100100011101110100000000101;
		b = 32'b00010111101001111001100100011100;
		correct = 32'b00110100101110110001110110100111;
		#400 //3.2179644e+17 * 1.0830772e-24 = 3.485304e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110001001010001110110001111;
		b = 32'b00011001110110110000100001101010;
		correct = 32'b00011000100011010100010110110111;
		#400 //0.16124557 * 2.2647468e-23 = 3.651804e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001111011100111000100101110100;
		b = 32'b00101001101111101010100011110010;
		correct = 32'b10111001101101010110000010111101;
		#400 //-4085871600.0 * 8.467002e-14 = -0.00034595086
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010110011111000110011111001101;
		b = 32'b11000001000010001010000111000110;
		correct = 32'b01011000000001101011011010100101;
		#400 //-69380688000000.0 * -8.539495 = 592476040000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001011101110101110001011111000;
		b = 32'b11111101001000110101001101111111;
		correct = 32'b11001001011011100111011011110000;
		#400 //7.19861e-32 * -1.3568606e+37 = -976751.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111111010000001010010010011010;
		b = 32'b00000101100001000001010001000101;
		correct = 32'b00000101010001101100100001000000;
		#400 //0.7525116 * 1.2420666e-35 = 9.3466954e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101010000110011110000111001000;
		b = 32'b11011011010010000010110110100011;
		correct = 32'b11000101111100001010011110100110;
		#400 //1.3667463e-13 * -5.6345173e+16 = -7700.956
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010001000010100011101100111100;
		b = 32'b01101100001011010000101010111011;
		correct = 32'b10111101101110101101111110100110;
		#400 //-1.0904533e-28 * 8.3677936e+26 = -0.09124689
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111101110100100010010110000010;
		b = 32'b10011100011100101110000111000001;
		correct = 32'b01011010110001110110000011000110;
		#400 //-3.491658e+37 * -8.0362863e-22 = 2.8059962e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010111011010011101110110010101;
		b = 32'b00001011001101011010000000111001;
		correct = 32'b10100011001001011110110000001001;
		#400 //-257137900000000.0 * 3.497987e-32 = -8.99465e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111000001010011110110110000001;
		b = 32'b10011010101010111010000010001000;
		correct = 32'b10010011011000111101100001101000;
		#400 //4.0513933e-05 * -7.0983295e-23 = -2.8758125e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100101110000110111110011100101;
		b = 32'b11000100111111001001101000011110;
		correct = 32'b11101011010000001110010010100001;
		#400 //1.1539567e+23 * -2020.8162 = -2.3319343e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011010110000011000110000000000;
		b = 32'b00110011001100010010110011000010;
		correct = 32'b00001110100001011111001110100011;
		#400 //8.004911e-23 * 4.125173e-08 = 3.3021645e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001010111110100001110101110100;
		b = 32'b11011001000011110000011010001100;
		correct = 32'b01100100100010111011110011011001;
		#400 //-8195770.0 * -2516132500000000.0 = 2.0621643e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111011111110100101111111111011;
		b = 32'b10001100101000101010100010001001;
		correct = 32'b00001001000111110001010110010010;
		#400 //-0.0076408363 * -2.5061485e-31 = 1.9149071e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101000100110010001001101110011;
		b = 32'b00110001000010101000101100001010;
		correct = 32'b01011010001001011010111100111111;
		#400 //5.783047e+24 * 2.0160678e-09 = 1.1659014e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100100111011110010101101011010;
		b = 32'b00101000011100111100011110101101;
		correct = 32'b10001101111000111100000010110011;
		#400 //-1.0372317e-16 * 1.35325075e-14 = -1.4036346e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111100010111100101100001100111;
		b = 32'b00000010100111101100010110110101;
		correct = 32'b00111111100010011110011001000111;
		#400 //4.6179317e+36 * 2.3329492e-37 = 1.07734
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011101000010010101111110110010;
		b = 32'b11000101001010100101001010010011;
		correct = 32'b01100010101101101100101110110111;
		#400 //-6.1867664e+17 * -2725.161 = 1.6859933e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011110001010000100010110100111;
		b = 32'b10000010011110101101001110011111;
		correct = 32'b10100001001001001101111100011111;
		#400 //3.0313203e+18 * -1.8427832e-37 = -5.586066e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111100001101110111001001011000;
		b = 32'b10011100011100000110100010111001;
		correct = 32'b11011001001011000100011000111110;
		#400 //3.810038e+36 * -7.954469e-22 = -3030683000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001000111100100000111100100111;
		b = 32'b00001101000100000010101110100110;
		correct = 32'b00010110100010000101000111001011;
		#400 //495737.22 * 4.4425966e-31 = 2.2023604e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110110000001111000011101011101;
		b = 32'b10011110100111100011001011011011;
		correct = 32'b01010101001001111000000011110000;
		#400 //-6.872125e+32 * -1.6749934e-20 = 11510764000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010000101011011101001000111;
		b = 32'b01111101100101110110110010000100;
		correct = 32'b11111000001100010010000010101111;
		#400 //-0.00057116564 * 2.515961e+37 = -1.4370304e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011101100010110000001010010;
		b = 32'b01001100001100011011011110110000;
		correct = 32'b11011000011101100100010110111101;
		#400 //-23249060.0 * 46587584.0 = -1083117540000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000110111111001000000010100011;
		b = 32'b00000111000100000100001100111100;
		correct = 32'b10001110100011100100101010101101;
		#400 //-32320.318 * 1.0853114e-34 = -3.5077613e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110110011101111100010111000111;
		b = 32'b00110011011101000110011111001101;
		correct = 32'b00101010011011001000110011111001;
		#400 //3.692099e-06 * 5.6905083e-08 = 2.100992e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101010101010001010011011010011;
		b = 32'b00011110001110101010001110011001;
		correct = 32'b11001001011101011110100111111001;
		#400 //-1.0194367e+26 * 9.880589e-21 = -1007263.56
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001111000001101011011100010111;
		b = 32'b01111010111011110111001000001010;
		correct = 32'b01001010011111000000000111100011;
		#400 //6.641972e-30 * 6.2163597e+35 = 4128888.8
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000101001100010001110100011000;
		b = 32'b01101011110011111010110000110100;
		correct = 32'b01110001100011111010110110101010;
		#400 //2833.8184 * 5.021217e+26 = 1.4229217e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011001011110101100110001000010;
		b = 32'b10111000000001010110111011011100;
		correct = 32'b00010010000000101011100010111010;
		#400 //-1.2965947e-23 * -3.1812917e-05 = 4.124846e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000110111100101010011101011;
		b = 32'b11110011010111110100100111011010;
		correct = 32'b01100100110000011110110000011100;
		#400 //-1.6176761e-09 * -1.7690736e+31 = 2.861788e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101110100101001010101011111110;
		b = 32'b10101011010001001100000010111100;
		correct = 32'b00011010011001001000010110110000;
		#400 //-6.760635e-11 * -6.990066e-13 = 4.7257287e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001100111110010001100000001111;
		b = 32'b11110011100110110011101001101100;
		correct = 32'b11000001000101110000101001101010;
		#400 //3.8379004e-31 * -2.4596892e+31 = -9.4400425
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111101100010001000011010011110;
		b = 32'b01011001001101111100000101101011;
		correct = 32'b01010111010000111111111011000011;
		#400 //0.06666301 * 3232661600000000.0 = 215498960000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110101101110110101000111000101;
		b = 32'b01001110100100100000001010000001;
		correct = 32'b01000100110101011010110011101111;
		#400 //1.3956384e-06 * 1224818800.0 = 1709.4042
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011011001101100011010011110000;
		b = 32'b00011100101110111010100111110001;
		correct = 32'b10111000100001011001000110100000;
		#400 //-5.128665e+16 * 1.2418551e-21 = -6.369059e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000101000000001000000111100010;
		b = 32'b10111011000011111011011011001011;
		correct = 32'b10000000100100000100100010011111;
		#400 //6.042387e-36 * -0.0021929021 = -1.3250363e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100011000100000110111000010100;
		b = 32'b00110111000100111111110111011011;
		correct = 32'b11011010101001101111110011011100;
		#400 //-2.664263e+21 * 8.820988e-06 = -2.3501434e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101100000111011001001111111011;
		b = 32'b00100010111001001111101010001000;
		correct = 32'b11001111100011001111001000000010;
		#400 //-7.620007e+26 * 6.2064784e-18 = -4729341000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111000100101011111110011001010;
		b = 32'b11000001000100010011110001010000;
		correct = 32'b00111010001010100010111100001001;
		#400 //-7.151959e-05 * -9.077225 = 0.0006491994
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110111011001000010111011111011;
		b = 32'b10100110011110001011111001110000;
		correct = 32'b10011110010111011011011101000010;
		#400 //1.36007975e-05 * -8.6300375e-16 = -1.17375394e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000100011010111001110011011100;
		b = 32'b10111111000110101111100000100010;
		correct = 32'b00000100000011101010000010111100;
		#400 //-2.7696144e-36 * -0.6053487 = 1.6765825e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011110001110110001101011010110;
		b = 32'b11010110111111010100111001101110;
		correct = 32'b01110101101110010010001011011000;
		#400 //-3.370581e+18 * -139256650000000.0 = 4.693758e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110110000110010001110101010100;
		b = 32'b01000111011010010000101111110101;
		correct = 32'b11111110000010110110001011011000;
		#400 //-7.763831e+32 * 59659.957 = -4.631898e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011011101011100100000011111111;
		b = 32'b11011111001000000110101010000111;
		correct = 32'b01111011010110100110001001000100;
		#400 //-9.809622e+16 * -1.15592e+19 = 1.1339138e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010100011010110101011100001001;
		b = 32'b11011101101011110000010101001100;
		correct = 32'b01110010101000001110010101011110;
		#400 //-4043110000000.0 * -1.5764462e+18 = 6.373746e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100011010011011001010100110110;
		b = 32'b11100111100001101101110111010110;
		correct = 32'b11001011010110001001110010000000;
		#400 //1.1144669e-17 * -1.2737785e+24 = -14195840.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100010010111000100010101100111;
		b = 32'b00011110100011010000010011110010;
		correct = 32'b10000001011100101010110011110110;
		#400 //-2.9852301e-18 * 1.4931001e-20 = -4.4572474e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000011001010111010111100000100;
		b = 32'b00000010011101110001100111110111;
		correct = 32'b10000110001001011011011101000111;
		#400 //-171.68365 * 1.8154146e-37 = -3.1167702e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011001011100100101100011111010;
		b = 32'b10010110101001110010011001011111;
		correct = 32'b00110000100111100011110001011110;
		#400 //-4263423400000000.0 * -2.700452e-25 = 1.151317e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011001011101010110101110010011;
		b = 32'b00111010111100101110101101101101;
		correct = 32'b11010100111010001110000101100011;
		#400 //-4317478000000000.0 * 0.0018533297 = -8001710000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010101101111000011010110011111;
		b = 32'b01001110110111110001111100101101;
		correct = 32'b01100101001001000000100110100001;
		#400 //25867310000000.0 * 1871681200.0 = 4.841536e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010101100100010001100010011100;
		b = 32'b10101111010001111110000000011000;
		correct = 32'b11000101011000101001001001001001;
		#400 //19941860000000.0 * -1.8178559e-10 = -3625.1428
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100100001101101110101010011100;
		b = 32'b11011001110101000010111100101101;
		correct = 32'b10111110100101111001101111111110;
		#400 //3.966368e-17 * -7465570700000000.0 = -0.296112
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111011011111110001100100100111;
		b = 32'b00111110111010100010011101111111;
		correct = 32'b00111010111010010101010001011001;
		#400 //0.0038924904 * 0.45733258 = 0.0017801627
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101100101111111100100010001101;
		b = 32'b01001101101100101101011010100101;
		correct = 32'b10111011000001011111101000111111;
		#400 //-5.450812e-12 * 375051420.0 = -0.0020443348
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000111101001110111010000101110;
		b = 32'b00110111000001001010000100000010;
		correct = 32'b10111111001011011000001001110010;
		#400 //-85736.36 * 7.905301e-06 = -0.6777717
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100110010010011101001111001001;
		b = 32'b11010011111010110000010100100011;
		correct = 32'b00111010101110010100100101110110;
		#400 //-7.0022906e-16 * -2018807000000.0 = 0.0014136273
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100010010100111111111010111101;
		b = 32'b10110110011100011001111111000100;
		correct = 32'b11011001010010000001011100011101;
		#400 //9.776547e+20 * -3.6004794e-06 = -3520025500000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011011011101010110001001111101;
		b = 32'b01000010100010011100100110010111;
		correct = 32'b00011110100001000001001011110000;
		#400 //2.0297748e-22 * 68.89373 = 1.3983876e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101010000101111100100010000111;
		b = 32'b00110001010100100100001011110101;
		correct = 32'b00011011111110010101010001100011;
		#400 //1.3481066e-13 * 3.0597083e-09 = 4.1248128e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111010001100001011100010011000;
		b = 32'b00101001111001110000001110010000;
		correct = 32'b11100100100111110111100100000111;
		#400 //-2.2939706e+35 * 1.0259079e-13 = -2.3534026e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000110101101010011101011101111;
		b = 32'b01110010100001110000110100010111;
		correct = 32'b11111001101111110011011010110001;
		#400 //-23197.467 * 5.3499265e+30 = -1.2410475e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010100011110011010111011010011;
		b = 32'b11111000111010011011000011000101;
		correct = 32'b01001101111000111110110010000110;
		#400 //-1.2605765e-26 * -3.7918453e+34 = 477991100.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000100010001011111111001100100;
		b = 32'b11001010111000001000000001110011;
		correct = 32'b10001111101011011010000111110000;
		#400 //2.327405e-36 * -7356473.5 = -1.7121493e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100101111100000100111000010111;
		b = 32'b00101101000101111111100000010000;
		correct = 32'b00010011100011101010011011101010;
		#400 //4.168628e-16 * 8.638437e-12 = 3.601043e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101010100100001111001111000011;
		b = 32'b01001110101011010011010000100101;
		correct = 32'b10111001110001000010010010000010;
		#400 //-2.5748682e-13 * 1452937900.0 = -0.00037411234
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010101100111101000000000100101;
		b = 32'b01100110011101001001000001010111;
		correct = 32'b00111100100101110110101110000001;
		#400 //6.401787e-26 * 2.8873e+23 = 0.018483879
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001011011101101011111001011011;
		b = 32'b01000111110101111001100101101111;
		correct = 32'b00010011110011111100110111000001;
		#400 //4.7521084e-32 * 110386.87 = 5.2457035e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111111001111100110110011000;
		b = 32'b01110010101001111011010001000100;
		correct = 32'b11101011000101111101101001011000;
		#400 //-2.7633083e-05 * 6.6434463e+30 = -1.835789e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011101011101111001110110110000;
		b = 32'b00010111111100001110111011001110;
		correct = 32'b10110101111010010000101011010001;
		#400 //-1.1151632e+18 * 1.5569919e-24 = -1.7363001e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011000011000111000010000000001;
		b = 32'b00110111111011110011100011010001;
		correct = 32'b01010000110101001001101010111100;
		#400 //1000624400000000.0 * 2.8517477e-05 = 28535284000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111110100001010000001111110100;
		b = 32'b10000100111000100001001010101100;
		correct = 32'b00000011111010101110111001100010;
		#400 //-0.25979578 * -5.3149492e-36 = 1.3808014e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100010000100001101011100011010;
		b = 32'b00101110001011110101100110010000;
		correct = 32'b10010000110001100110101101101110;
		#400 //-1.9629513e-18 * 3.986994e-11 = -7.826275e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011100011000110101111000000100;
		b = 32'b10101010010010000001011011100000;
		correct = 32'b01000111001100011011010111000100;
		#400 //-2.5599276e+17 * -1.7771505e-13 = 45493.766
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101110110011111100010000000101;
		b = 32'b01101011000010011001000111101111;
		correct = 32'b01011010010111110100110010101101;
		#400 //9.44809e-11 * 1.6631199e+26 = 1.5713306e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011100101000011111100100100100;
		b = 32'b11001001100011111000101111001010;
		correct = 32'b01100110101101011010010100111010;
		#400 //-3.6473123e+17 * -1175929.2 = 4.288981e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010101111110011011101000000;
		b = 32'b11000110010111100111111000100000;
		correct = 32'b01000001101001100011000000011111;
		#400 //-0.0014588609 * -14239.531 = 20.773497
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101111100001110011001100111011;
		b = 32'b01001100000001010011000101000011;
		correct = 32'b10111100000011001010111101000100;
		#400 //-2.4592758e-10 * 34915596.0 = -0.008586708
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001001101101000000000110101110;
		b = 32'b01101011000000100000111110110001;
		correct = 32'b11110101001101101110011111000110;
		#400 //-1474613.8 * 1.5723446e+26 = -2.318601e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110100010001001111010101101111;
		b = 32'b10100001010001000011110011101010;
		correct = 32'b01010110000101101111101011000111;
		#400 //-6.241871e+31 * -6.6488e-19 = 41500956000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010110010110101001100001110111;
		b = 32'b11100010000100010011010010100000;
		correct = 32'b11111000111101111111101010010110;
		#400 //60087090000000.0 * -6.696425e+20 = -4.023687e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111010001011100100000001000000;
		b = 32'b10101001011011111100111111000111;
		correct = 32'b11100100001000110011101101101001;
		#400 //2.261907e+35 * -5.324888e-14 = -1.2044401e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110110011111011011110110111100;
		b = 32'b01100011111111101011011110011100;
		correct = 32'b01011010111111000111100000111110;
		#400 //3.7810378e-06 * 9.397407e+21 = 3.553195e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110000010110010101000110000101;
		b = 32'b01100111111001110110011101111010;
		correct = 32'b01011000110001000111000001100110;
		#400 //7.9059986e-10 * 2.1855509e+24 = 1727896200000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111010011000000111101100010100;
		b = 32'b10101011000010010010011100110101;
		correct = 32'b01100101111100001000100001111110;
		#400 //-2.913927e+35 * -4.872659e-13 = 1.4198572e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010101011010111100001111110111;
		b = 32'b01010010010000111001111011011110;
		correct = 32'b11101000001101000010100010010101;
		#400 //-16201681000000.0 * 210046000000.0 = -3.4030983e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010101010000011100100100101100;
		b = 32'b01100100010100101111010110100001;
		correct = 32'b11111010000111111011000011110101;
		#400 //-13316861000000.0 * 1.5566063e+22 = -2.0729108e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100001101000011100111001011000;
		b = 32'b10110100111110111101110100011011;
		correct = 32'b11010111000111110011000100010000;
		#400 //3.730993e+20 * -4.691327e-07 = -175033070000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000000010111111001001111101111;
		b = 32'b00000001011111011110000111111100;
		correct = 32'b00000010010111011011101010010000;
		#400 //3.4934042 * 4.6630897e-38 = 1.6290057e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011001001001110011000101000011;
		b = 32'b11001110101010100111110110100001;
		correct = 32'b11101000010111101011000110000101;
		#400 //2941280300000000.0 * -1430180000.0 = -4.20656e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011100110000110000010100110111;
		b = 32'b00101000001110111110010100110111;
		correct = 32'b11000101100011110010001101101101;
		#400 //-4.3914683e+17 * 1.0430288e-14 = -4580.428
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101101010001000010011011011011;
		b = 32'b10001011000000011110100001010101;
		correct = 32'b10111000110001110001001100110001;
		#400 //3.7941272e+27 * -2.5019283e-32 = -9.492634e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101111010110111011101011111110;
		b = 32'b00101001101010110101000001100111;
		correct = 32'b00011001100100110000101011101011;
		#400 //1.9984367e-10 * 7.607873e-14 = 1.5203853e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110011100000100010000011101100;
		b = 32'b00111110111101101001010000011001;
		correct = 32'b00110010111110101010110111010101;
		#400 //6.059585e-08 * 0.48159865 = 2.918288e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001000001100001001010000111111;
		b = 32'b01100110101010101110100001000001;
		correct = 32'b11101111011010111100010101001010;
		#400 //-180816.98 * 4.035433e+23 = -7.2967485e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000011100100101010111111101101;
		b = 32'b11010010000010100010001011110000;
		correct = 32'b10010110000111100100110110110101;
		#400 //8.621499e-37 * -148322910000.0 = -1.2787658e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011111001010010001110011001111;
		b = 32'b11010010100000111000111001110100;
		correct = 32'b01110010001011011100111110110001;
		#400 //-1.2185842e+19 * -282515340000.0 = 3.4426874e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111000010010001100111000101100;
		b = 32'b10111101001010001011011110101011;
		correct = 32'b11110110000001000101011101011110;
		#400 //1.6291266e+34 * -0.041190784 = -6.7105e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110111111011011011100110100111;
		b = 32'b01000000001100001111010000011100;
		correct = 32'b11111000101001000101001001010010;
		#400 //-9.64328e+33 * 2.7648993 = -2.6662698e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100111101110100011011001110;
		b = 32'b10100010000001011111101000100011;
		correct = 32'b10100111100000010110100101100110;
		#400 //1978.2126 * -1.8157282e-18 = -3.5918966e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011111011110011101110100101101;
		b = 32'b01000100111010011001001001001011;
		correct = 32'b00100100111000111111100100010111;
		#400 //5.2910753e-20 * 1868.5717 = 9.886753e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110010100110001010001110000010;
		b = 32'b01111111011100000110111111011100;
		correct = 32'b01110010100011110101101111111100;
		#400 //1.7769484e-08 * 3.1959553e+38 = 5.6790475e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101111001111100110100010010110;
		b = 32'b00000101000000001000101111100011;
		correct = 32'b00110100101111110011100010101101;
		#400 //5.892859e+28 * 6.044224e-36 = 3.561776e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101101110000011001001111101001;
		b = 32'b11000001110010110011010001000101;
		correct = 32'b01110000000110011010011111010000;
		#400 //-7.4886774e+27 * -25.400522 = 1.9021632e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001111111101010010010110110101;
		b = 32'b10001100111000110111100000110110;
		correct = 32'b00011101010110011101001110001101;
		#400 //-8225778000.0 * -3.5047237e-31 = 2.882908e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011110110010011110101010001001;
		b = 32'b11011011101010010101000101110110;
		correct = 32'b11111011000001011000110000010101;
		#400 //7.274796e+18 * -9.531768e+16 = -6.934167e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110010111011101011111111011100;
		b = 32'b00011001100001111110110011000100;
		correct = 32'b01001100111111011000011111111001;
		#400 //9.45784e+30 * 1.4054302e-23 = 132923336.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101010111011101000010010100101;
		b = 32'b10011001001011010000100110111110;
		correct = 32'b01000100101000010011100010110111;
		#400 //-1.4417537e+26 * -8.945858e-24 = 1289.7723
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011011110000100110000001011111;
		b = 32'b10110110010110101100011100100000;
		correct = 32'b11010010101001100001110101000010;
		#400 //1.0942421e+17 * -3.2600437e-06 = -356727720000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110110010110111111001101110011;
		b = 32'b01000010010000111010001000010011;
		correct = 32'b11111001001010000001010110110001;
		#400 //-1.1152839e+33 * 48.908276 = -5.4546614e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011101010000000000111010001000;
		b = 32'b11011101101000111110101001010100;
		correct = 32'b10111011011101011111001000011010;
		#400 //2.54185e-21 * -1.4764182e+18 = -0.0037528337
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110001101111110111110100010001;
		b = 32'b01010000011111101111100000111101;
		correct = 32'b11000010101111101011011111000110;
		#400 //-5.57305e-09 * 17110726000.0 = -95.35893
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010000010110001010010000000001;
		b = 32'b00001111110010000110111101101000;
		correct = 32'b00100000101010011001111001101000;
		#400 //14538507000.0 * 1.9764435e-29 = 2.8734538e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101000110010101010001101000111;
		b = 32'b00100110110001100010010111101010;
		correct = 32'b10010000000111001101100001001100;
		#400 //-2.2497315e-14 * 1.3749287e-15 = -3.0932204e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001111001000000110011011111100;
		b = 32'b10110010001001101000111011100000;
		correct = 32'b10000001110100001011100010011010;
		#400 //7.908443e-30 * -9.694958e-09 = -7.6672023e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010000101000110100000101101101;
		b = 32'b11010110101110010101110000011011;
		correct = 32'b10100111111011000110101000001001;
		#400 //6.439297e-29 * -101902620000000.0 = -6.561812e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010101101010101011011111100111;
		b = 32'b00110000000001111110011100001110;
		correct = 32'b00000110001101010100001000100000;
		#400 //6.89526e-26 * 4.944106e-10 = 3.4090897e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111001001001001110100110000;
		b = 32'b01101010011101000001100010001000;
		correct = 32'b01110010000111001111010110011000;
		#400 //42141.188 * 7.3773436e+25 = 3.1089002e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110110101000010100001010001000;
		b = 32'b00111010100101101011010001010101;
		correct = 32'b01110001101111011101110100101000;
		#400 //1.6353695e+33 * 0.0011497835 = 1.8803209e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001001101001011100000010101111;
		b = 32'b11101000111100011111000101000101;
		correct = 32'b01110011000111001010011010011100;
		#400 //-1357845.9 * -9.1403277e+24 = 1.2411156e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001101010100011001011111110010;
		b = 32'b11100111011011001101101101010110;
		correct = 32'b00110101010000011110101110100110;
		#400 //-6.4585995e-31 * -1.1185245e+24 = 7.2241016e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101011001010101000101100111110;
		b = 32'b11110001001001110001100001001101;
		correct = 32'b11011100110111101010001000001100;
		#400 //6.058937e-13 * -8.27414e+29 = -5.0132494e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001101001110101100000011101011;
		b = 32'b11110001100010000010110101011110;
		correct = 32'b11111111010001101010111100101011;
		#400 //195825330.0 * -1.3486338e+30 = -2.6409667e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011010101101011000001010101110;
		b = 32'b01101101101000111101010101110110;
		correct = 32'b01001000111010000101001100011100;
		#400 //7.507097e-23 * 6.3380144e+27 = 475800.88
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010110100010000101111011011101;
		b = 32'b10000010000001010000010110011001;
		correct = 32'b10011001000011011011100010001000;
		#400 //74970510000000.0 * -9.772903e-38 = -7.326795e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100100001000001010011100011010;
		b = 32'b10001111100101010100100101011111;
		correct = 32'b00110100001110110101111010011011;
		#400 //-1.185408e+22 * -1.4720796e-29 = 1.745015e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110001100111100010111010100101;
		b = 32'b00010010011011000010101001111000;
		correct = 32'b01000100100100011110110100111110;
		#400 //1.5665607e+30 * 7.4520816e-28 = 1167.4138
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000100101100010010100001001110;
		b = 32'b01101111100000100011001011111111;
		correct = 32'b11110100101101000011001110000100;
		#400 //-1417.2595 * 8.05894e+28 = -1.142161e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011000011000111101001011000110;
		b = 32'b10100100101101010111001001000010;
		correct = 32'b10111101101000010111100110110101;
		#400 //1001977600000000.0 * -7.86898e-17 = -0.07884542
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010111000110100011011110110;
		b = 32'b10101011001101101111111110010100;
		correct = 32'b00100110101000100111011101011010;
		#400 //-0.0017339874 * -6.5014075e-13 = 1.1273358e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000000100100010110101100100110;
		b = 32'b01000101111000111100001011100001;
		correct = 32'b10000111000000010110000010110110;
		#400 //-1.3354585e-38 * 7288.36 = -9.733302e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101100101111100000000011001111;
		b = 32'b01000001000000101011011001101011;
		correct = 32'b00101110010000100000011110011010;
		#400 //5.4002146e-12 * 8.169536 = 4.4117245e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101110000001000010101100110111;
		b = 32'b10110010110110111010000001000000;
		correct = 32'b10100001011000101100011101101000;
		#400 //3.0051708e-11 * -2.5567829e-08 = -7.683569e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100010010010001111011110101010;
		b = 32'b10001010100011101001010100100011;
		correct = 32'b10101101010111111101110011101000;
		#400 //9.267987e+20 * -1.3730202e-32 = -1.27251334e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011111101000100011011000100101;
		b = 32'b11110001010011100110110010101101;
		correct = 32'b11010001100000101100110001101110;
		#400 //6.8699243e-20 * -1.0221647e+30 = -70221940000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111110011000101011100010010;
		b = 32'b10100011110000001000011010000001;
		correct = 32'b10101100000110011010110010101010;
		#400 //104622.14 * -2.0873646e-17 = -2.1838456e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011100100000110000001011000011;
		b = 32'b10101001010010101010111001001111;
		correct = 32'b01000110010011110111001011000100;
		#400 //-2.9501007e+17 * -4.50042e-14 = 13276.691
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001110001110000000111000111010;
		b = 32'b10000110101000010110000100000101;
		correct = 32'b10010101011010000000110101100111;
		#400 //771985000.0 * -6.0704026e-35 = -4.68626e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100100111011100110100101011101;
		b = 32'b10101011011101011001110110000111;
		correct = 32'b01010000111001001011110110001010;
		#400 //-3.5183339e+22 * -8.72601e-13 = 30701015000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101010101010110000000100101011;
		b = 32'b01011100000011001010101001010101;
		correct = 32'b11000111001110111110110011010110;
		#400 //-3.0376512e-13 * 1.5837512e+17 = -48108.836
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010011111101100111100111000000;
		b = 32'b00110101001111101001011011010011;
		correct = 32'b00001001101101110111111110010011;
		#400 //6.2219185e-27 * 7.0999994e-07 = 4.4175618e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100001110100011011111011111;
		b = 32'b01010100110101101110001110001110;
		correct = 32'b01011001100111000101000000111011;
		#400 //744.873 * 7383526000000.0 = 5499789000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100110110000001010000101110010;
		b = 32'b11110110100100010110000010110010;
		correct = 32'b11011101110110101100100001101000;
		#400 //1.3366436e-15 * -1.4743052e+33 = -1.9706206e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100100110011010011011001011001;
		b = 32'b01101100010101110100101100011000;
		correct = 32'b01010001101011001001010011010111;
		#400 //8.8996647e-17 * 1.0410947e+27 = 92653940000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010000011110011010010101100110;
		b = 32'b01010110101000100111101100000011;
		correct = 32'b10100111100111100111001010100000;
		#400 //-4.923401e-29 * 89324610000000.0 = -4.3978086e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111010011001110110001000111100;
		b = 32'b01111111010011001000010111010000;
		correct = 32'b01111010001110001101101100111010;
		#400 //0.0008826589 * 2.718573e+38 = 2.3995727e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110000001101100101100001101000;
		b = 32'b01010101011100011010101001001100;
		correct = 32'b01000110001011000010001010000111;
		#400 //6.6336847e-10 * 16607108000000.0 = 11016.632
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101100011011000110000000010000;
		b = 32'b00110001111011000110100000000100;
		correct = 32'b00011110110110100100100010011001;
		#400 //3.3590943e-12 * 6.880329e-09 = 2.3111673e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010111010000011001001001100100;
		b = 32'b10101100111011001001101010011101;
		correct = 32'b01000100101100101110011111011101;
		#400 //-212834490000000.0 * -6.724689e-12 = 1431.2457
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000010101001010100011001000001;
		b = 32'b00100011010101101000011011010011;
		correct = 32'b10100110100010100111111111000101;
		#400 //-82.637215 * 1.1629513e-17 = -9.610306e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111011000110010110110110011110;
		b = 32'b00001100000111110010101110000011;
		correct = 32'b00000111101111101100101001010010;
		#400 //0.0023411284 * 1.2262008e-31 = 2.8706936e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101001101111001001101010110011;
		b = 32'b00001010011010001011010101010111;
		correct = 32'b00110100101010110111000111001100;
		#400 //2.8501075e+25 * 1.12045e-32 = 3.193403e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111101111110010001010011000100;
		b = 32'b10100011001001111101011011010101;
		correct = 32'b11100001101000110100110110010010;
		#400 //4.13857e+37 * -9.098581e-18 = -3.765511e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000000111000110111110000111110;
		b = 32'b01001001110101100100011110111001;
		correct = 32'b01001011001111100110100110011000;
		#400 //7.1089163 * 1755383.1 = 12478872.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000111101011000111101111110111;
		b = 32'b01010100000000011100011111011111;
		correct = 32'b11011100001011101110001001000100;
		#400 //-88311.93 * 2229616200000.0 = -1.9690171e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100101101100111000110001101100;
		b = 32'b01010100001111110101000011011100;
		correct = 32'b01111010100001100010111001111011;
		#400 //1.0598674e+23 * 3286781400000.0 = 3.4835526e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001011001000010010001111110000;
		b = 32'b00111010101101011100001000110011;
		correct = 32'b01000110011001001101000101001100;
		#400 //10560496.0 * 0.001386708 = 14644.324
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100100100100010111011010101011;
		b = 32'b00100010111111011110110000100011;
		correct = 32'b10001000000100000100100001110100;
		#400 //-6.308476e-17 * 6.8825807e-18 = -4.341859e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101011100011101011010110111011;
		b = 32'b11101101010000010101101100010010;
		correct = 32'b11011001010101111001001110001101;
		#400 //1.0140147e-12 * -3.740044e+27 = -3792459600000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101110000100111111011010000001;
		b = 32'b01001111011110000110011001001100;
		correct = 32'b10111110000011111001000111101101;
		#400 //-3.364287e-11 * 4167453700.0 = -0.1402051
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011011101000111001101010110000;
		b = 32'b01010101101000100010111110001011;
		correct = 32'b01110001110011110100110010001011;
		#400 //9.2101e+16 * 22290635000000.0 = 2.0529898e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001000011110101011101110111001;
		b = 32'b00100111011011010000000000000100;
		correct = 32'b10110000011010000001111111001110;
		#400 //-256750.89 * 3.2890366e-15 = -8.4446306e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100100000010011111110001111;
		b = 32'b01010010011101001111000111111111;
		correct = 32'b01010111011101110101010110000100;
		#400 //1033.9862 * 263008010000.0 = 271946660000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010111000000010001011010000110;
		b = 32'b11001101101010010001000010111111;
		correct = 32'b10100101001010101000000010100000;
		#400 //4.1710577e-25 * -354555870.0 = -1.478873e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000101111111110111000101100000;
		b = 32'b01000111100110100111011110011110;
		correct = 32'b01001110000110100010000110001111;
		#400 //8174.172 * 79087.234 = 646472640.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101011111110001000101011101011;
		b = 32'b01010000010101010001101000100001;
		correct = 32'b00111100110011101110010011110100;
		#400 //1.7660017e-12 * 14301038000.0 = 0.025255658
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101100010100100110110010010000;
		b = 32'b00011100111101001001010000010011;
		correct = 32'b01001001110010010000100100110000;
		#400 //1.0175484e+27 * 1.6184842e-21 = 1646886.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111000110000001011101000110000;
		b = 32'b10100110010010110010101001100111;
		correct = 32'b00011111100110001111001110010000;
		#400 //-9.1899536e-05 * -7.048724e-16 = 6.4777444e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111111101000011101001011001010;
		b = 32'b01111000111010110011010101111001;
		correct = 32'b01111001000101001010111001001101;
		#400 //1.2642453 * 3.8164822e+34 = 4.82497e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111011000101101000000000010;
		b = 32'b10001000101111100000010110100011;
		correct = 32'b00000000101010000101101101100000;
		#400 //-1.351908e-05 * -1.1436534e-33 = 1.5461143e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011110001110111100011000000111;
		b = 32'b11001110100001011010010010111001;
		correct = 32'b01101101010001000000110101101000;
		#400 //-3.3826275e+18 * -1121082500.0 = 3.7922043e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001001000100011010001001110011;
		b = 32'b11001000011101110111000000000101;
		correct = 32'b01010010000011001100001101110111;
		#400 //-596519.2 * -253376.08 = 151143700000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000000110101001000110001010;
		b = 32'b11000100010111100110101011011001;
		correct = 32'b00110101000001100100101010111001;
		#400 //-5.6231697e-10 * -889.6695 = 5.0027626e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100010101100101101110111100101;
		b = 32'b00010011100011011100011110010001;
		correct = 32'b10110110110001100001111101001110;
		#400 //-1.6497548e+21 * 3.579019e-27 = -5.904504e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010111010111111011110001111011;
		b = 32'b01100101010101001110101001100111;
		correct = 32'b11111101001110100001010011110010;
		#400 //-246000610000000.0 * 6.2841603e+22 = -1.5459073e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100111001010101101000101101001;
		b = 32'b11110111111011010011000110101110;
		correct = 32'b01011111100111100100010100000100;
		#400 //-2.370576e-15 * -9.621734e+33 = 2.2809052e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000010110010010000001010111101;
		b = 32'b11100011111010011000100010111010;
		correct = 32'b11100111001101110101111011011010;
		#400 //100.50535 * -8.615887e+21 = -8.659428e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111100000001010100001000001010;
		b = 32'b11011000101000010011101101000011;
		correct = 32'b01010101001001111101101011000011;
		#400 //-0.008133421 * -1418207200000000.0 = 11534876000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110011000111100001001001011101;
		b = 32'b10010100011110110100010100001011;
		correct = 32'b11001000000110110010011010100011;
		#400 //1.2523733e+31 * -1.2685878e-26 = -158874.55
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111000000111011100011111010100;
		b = 32'b10011010000001001000110110100110;
		correct = 32'b11010010101000110110010010101101;
		#400 //1.2800681e+34 * -2.7411383e-23 = -350884360000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001001111110100000101100100111;
		b = 32'b10000110111110010010101111001101;
		correct = 32'b00010001011100110101111110100001;
		#400 //-2048356.9 * -9.372775e-35 = 1.9198788e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011010001010000101101101011011;
		b = 32'b10100000101010010111111101111000;
		correct = 32'b10111011010111101111000001000111;
		#400 //1.1847061e+16 * -2.8714065e-19 = -0.0034017728
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111001111001101000000011101100;
		b = 32'b00111111101010100101010101001101;
		correct = 32'b10111010000110010101111001101011;
		#400 //-0.00043965073 * 1.3307282 = -0.0005850556
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011000100100101100001011101000;
		b = 32'b01111010010100011110111110111101;
		correct = 32'b01010011011100001011010100011111;
		#400 //3.793692e-24 * 2.7251313e+35 = 1033830860000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011111011010000000101101101100;
		b = 32'b00111111000101010000011101011010;
		correct = 32'b01011111000001110001010101010000;
		#400 //1.6720577e+19 * 0.5821434 = 9.733774e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101010001100000011000010000010;
		b = 32'b00111110000000001001101001110001;
		correct = 32'b01101000101100010000010100011000;
		#400 //5.3250004e+25 * 0.12558915 = 6.6876226e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100110010110001100100111011010;
		b = 32'b11001001011010010110011111101101;
		correct = 32'b01110000010001011010011110111001;
		#400 //-2.5593867e+23 * -956030.8 = 2.4468524e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011111101110111000111100010000;
		b = 32'b00101100111110111101110100100001;
		correct = 32'b01001101001110001000011101000111;
		#400 //2.7030077e+19 * 7.1583993e-12 = 193492080.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001111011001101010011011010111;
		b = 32'b00111101100010111111000101010011;
		correct = 32'b00001101011111000010110000001001;
		#400 //1.1372008e-29 * 0.06833138 = 7.77065e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010000110111111101000101001110;
		b = 32'b11101011110111000111100101101011;
		correct = 32'b11111101010000001100001000000111;
		#400 //30040290000.0 * -5.3307412e+26 = -1.6013701e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010110100110010111001110001010;
		b = 32'b00110000010111110101011000111101;
		correct = 32'b01000111100001011101111101010111;
		#400 //84360760000000.0 * 8.124948e-10 = 68542.68
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110100011100001010111001111100;
		b = 32'b10101010000100100111001101100110;
		correct = 32'b11011111000010011011000000000001;
		#400 //7.6275037e+31 * -1.3007442e-13 = -9.921431e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001010111000111001011000001101;
		b = 32'b01101100011011100110100010010111;
		correct = 32'b11110111110100111111001001111011;
		#400 //-7457542.5 * 1.152873e+27 = -8.5975994e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001010000011000001010100000110;
		b = 32'b11001010110000110111100100111010;
		correct = 32'b00010101010101011110110010110010;
		#400 //-6.744709e-33 * -6405277.0 = 4.3201727e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111000111010011000101000100010;
		b = 32'b10011101101101101100111001101001;
		correct = 32'b01010111001001101100010010000001;
		#400 //-3.7893964e+34 * -4.838842e-21 = 183362900000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110110000100010000111001111010;
		b = 32'b01000001000101001010011111011010;
		correct = 32'b00110111101010000111011011110101;
		#400 //2.161511e-06 * 9.290979 = 2.0082554e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011001110011000000011011101101;
		b = 32'b11111110001000110111110100011011;
		correct = 32'b11011000100000100100110000011110;
		#400 //2.1095903e-23 * -5.4328437e+37 = -1146107500000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000000001011011110001011110011;
		b = 32'b01101100010101001010010100011110;
		correct = 32'b01101101000100000111000000011001;
		#400 //2.716977 * 1.0282881e+27 = 2.793835e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101011111010010110100001110000;
		b = 32'b01001001101100110100010100011011;
		correct = 32'b01110110001000110111001100001000;
		#400 //5.643458e+26 * 1468579.4 = 8.287866e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001111101110001011001011101100;
		b = 32'b01010110101001001010011111000001;
		correct = 32'b10100110111011011001011101001110;
		#400 //-1.8212719e-29 * 90520200000000.0 = -1.648619e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001010010111101010000010000110;
		b = 32'b11001000100000010110100100100110;
		correct = 32'b10010011011000010001010010101001;
		#400 //1.0719102e-32 * -265033.2 = -2.8409179e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000111000001100001000010001001;
		b = 32'b01110001001001100110010000000111;
		correct = 32'b00111000101011100100011000110110;
		#400 //1.0085899e-34 * 8.23927e+29 = 8.310044e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100100010111100110010111110001;
		b = 32'b11010000111111010110001101000001;
		correct = 32'b10110101110111000010000011111001;
		#400 //4.8224924e-17 * -34009123000.0 = -1.6400874e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111110110000110001111100100100;
		b = 32'b00100000111111001001110010001110;
		correct = 32'b10100000010000001000100111111011;
		#400 //-0.38109696 * 4.279406e-19 = -1.6308686e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110111110011011011111000000000;
		b = 32'b01111110000001001001010001000101;
		correct = 32'b01110110010101010001101001000011;
		#400 //2.452638e-05 * 4.405699e+37 = 1.0805585e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101111101011110001100101110010;
		b = 32'b00101010101000101110010011010111;
		correct = 32'b00011010110111101101010101000000;
		#400 //3.1850395e-10 * 2.893577e-13 = 9.216157e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100100110001110010011001101001;
		b = 32'b01110011010111010101001010100000;
		correct = 32'b11011000101011000010110001101111;
		#400 //-8.636756e-17 * 1.7534995e+31 = -1514454700000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111100011110100101111001100001;
		b = 32'b11100111111010110000100100100010;
		correct = 32'b11100100111001011101110110010010;
		#400 //0.015281291 * -2.2198492e+24 = -3.3922162e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010010110010000101101111011110;
		b = 32'b10111010101000101110011111010111;
		correct = 32'b10001101111111101111111100101011;
		#400 //1.26444215e-27 * -0.0012428713 = -1.5715388e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010010001101100001111010011100;
		b = 32'b01100011011110001111110001001111;
		correct = 32'b00110110001100010010000100100101;
		#400 //5.7466803e-28 * 4.5929733e+21 = 2.6394348e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111011100100000010100001101010;
		b = 32'b10111101110001110000111101111010;
		correct = 32'b01111001111000000011000001000011;
		#400 //-1.4970209e+36 * -0.09719749 = 1.4550667e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001100110000000110110100111111;
		b = 32'b10011100000100000001011100100100;
		correct = 32'b00101001010110001001110110110001;
		#400 //-100887030.0 * -4.767551e-22 = 4.809841e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101001011100110100010000010000;
		b = 32'b11000001101100011111101010101111;
		correct = 32'b11101011101010010010000001000110;
		#400 //1.8380649e+25 * -22.247404 = -4.0892174e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101111111001100111010011000100;
		b = 32'b01110011110010000011011001111100;
		correct = 32'b11100100001101000011110001000101;
		#400 //-4.1919723e-10 * 3.172499e+31 = -1.3299027e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011001011011111100010111111101;
		b = 32'b01010110111100101100110000101011;
		correct = 32'b10110000111000110110100001100011;
		#400 //-1.2395994e-23 * 133479354000000.0 = -1.6546092e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110110001110100010000110001100;
		b = 32'b00111000111000101111110010011110;
		correct = 32'b11101111101001010000100101001001;
		#400 //-9.437965e+32 * 0.000108235734 = -1.021525e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011011110110011100111111111101;
		b = 32'b00101101000001001111000001111110;
		correct = 32'b01001001011000100011011110111001;
		#400 //1.2261751e+17 * 7.556731e-12 = 926587.56
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110000010010001001101100111110;
		b = 32'b10111111001000100010100101001101;
		correct = 32'b01101111111111100010010100110101;
		#400 //-2.4833871e+29 * -0.6334427 = 1.5730835e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011101010001011001001010111000;
		b = 32'b10110111000000001000001101000111;
		correct = 32'b00010100110001100101110101011010;
		#400 //-2.6148585e-21 * -7.65996e-06 = 2.0029711e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100000011000011001010001110111;
		b = 32'b00100101011111011101010000111010;
		correct = 32'b10000110010111111010101010111100;
		#400 //-1.9107364e-19 * 2.2016157e-16 = -4.2067074e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101110100100000111010010111110;
		b = 32'b00101101001100110110101101000000;
		correct = 32'b01011100010010100111110001001100;
		#400 //2.2353487e+28 * 1.0198786e-11 = 2.2797844e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010100000110110011100011001;
		b = 32'b11011001010110010000001100111101;
		correct = 32'b01010100010111101100100000011011;
		#400 //-0.0010025232 * -3817727000000000.0 = 3827359800000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010111001010110100101010010011;
		b = 32'b10001100010101101110110011000101;
		correct = 32'b10100100000011111100111011000011;
		#400 //188336780000000.0 * -1.655721e-31 = -3.1183316e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010001101011011110110101100000;
		b = 32'b01000010011011011100010111101100;
		correct = 32'b01010100101000011000101100111010;
		#400 //93376480000.0 * 59.443283 = 5550604600000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111111010110100111000111000000;
		b = 32'b10001000100101011001001101010110;
		correct = 32'b10001000011111110100001111011011;
		#400 //0.8532982 * -9.00225e-34 = -7.6816035e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000010000010011011111001010101;
		b = 32'b11101001110110011011011101000001;
		correct = 32'b10101100011010100100100111100000;
		#400 //1.0119793e-37 * -3.2900287e+25 = -3.3294409e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001100111111000000000100010101;
		b = 32'b11011001110111000100110101110100;
		correct = 32'b10100111010110001101110100101101;
		#400 //3.88274e-31 * -7751207000000000.0 = -3.0095921e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000101110111100001101010010111;
		b = 32'b00111010111010101110011000101000;
		correct = 32'b01000001010010111100101111111101;
		#400 //7107.3237 * 0.0017921375 = 12.737302
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110001011110110000000001010111;
		b = 32'b00111011100000100110011001010010;
		correct = 32'b00101101011111111011010011111101;
		#400 //3.65255e-09 * 0.0039794827 = 1.4535259e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101000011001111100000110100001;
		b = 32'b00111100000000111110100100110001;
		correct = 32'b00100100111011101101011001100010;
		#400 //1.28650625e-14 * 0.008051203 = 1.03579225e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010010100000111111110001111100;
		b = 32'b11111110010010011010001111010001;
		correct = 32'b01010001010011111110101101100110;
		#400 //-8.3295045e-28 * -6.7006353e+37 = 55812973000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010101011010001000000010111101;
		b = 32'b10110110101000010001110110010110;
		correct = 32'b11001100100100100101001111010110;
		#400 //15977477000000.0 * -4.801618e-06 = -76717740.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110111110010100100001011111001;
		b = 32'b00101101101111001001000110110001;
		correct = 32'b01100110000101001111110001001011;
		#400 //8.204706e+33 * 2.1437825e-11 = 1.7589106e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101111000010001111010111101001;
		b = 32'b10010110100000010000101110111011;
		correct = 32'b10000110000010100001010001100010;
		#400 //1.2456493e-10 * -2.0848477e-25 = -2.596989e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111100101110000111011111011001;
		b = 32'b01110110111111000001110011010100;
		correct = 32'b11110100001101011010101010111111;
		#400 //-0.022518085 * 2.5567256e+33 = -5.7572563e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111110010111110101010110110010;
		b = 32'b01000011000011010011010101011100;
		correct = 32'b11000001111101100110000110000000;
		#400 //-0.21810034 * 141.20844 = -30.797607
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000110111100010111101000111001;
		b = 32'b10010000101100100001100010000011;
		correct = 32'b00011000001001111111111000011011;
		#400 //-30909.111 * -7.0246387e-29 = 2.1712535e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111001001001101011100100001;
		b = 32'b01101100001010111001000110000011;
		correct = 32'b11100011110111001111001011001010;
		#400 //-9.82525e-06 * 8.296539e+26 = -8.151557e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011010010100110001010110100100;
		b = 32'b01010110000000011000011100001010;
		correct = 32'b10110000110101011001101010000001;
		#400 //-4.365126e-23 * 35604247000000.0 = -1.5541702e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111010010010010100111011010100;
		b = 32'b01100110011010000011010100011001;
		correct = 32'b01100001001101101001100100110001;
		#400 //0.0007679288 * 2.7414213e+23 = 2.1052163e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000100011111011000100000111110;
		b = 32'b00011100111010011010010100011100;
		correct = 32'b10100001111001110110010010000101;
		#400 //-1014.1288 * 1.5461326e-21 = -1.5679776e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000110111001110111110011100000;
		b = 32'b11101101010010011111100011101010;
		correct = 32'b00110100101101101010001000100000;
		#400 //-8.707603e-35 * -3.9067129e+27 = 3.4018103e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100110110001110101011100001101;
		b = 32'b11001110101010000011111011011101;
		correct = 32'b01110110000000110000001000010100;
		#400 //-4.7067837e+23 * -1411346000.0 = 6.642901e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101101100110110101010100000001;
		b = 32'b11001111010000110101100000010001;
		correct = 32'b01111101011011010000111001011111;
		#400 //-6.0091175e+27 * -3277328600.0 = 1.9693853e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011100001001111110000111010010;
		b = 32'b11010011111001100101000100100000;
		correct = 32'b10110000100101110000101000010110;
		#400 //5.554753e-22 * -1978407000000.0 = -1.0989563e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111010111011101010011001110011;
		b = 32'b01011111100100111111011001111001;
		correct = 32'b01011011000010011110111101011001;
		#400 //0.0018207565 * 2.1323684e+19 = 3.8825237e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100011000011110100110011001000;
		b = 32'b11000000110011101110001011001110;
		correct = 32'b00100100011001111001110101111100;
		#400 //-7.768305e-18 * -6.465186 = 5.0223535e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111100011111011001011000011100;
		b = 32'b10010110100001110100010011100110;
		correct = 32'b01010011100001011111111001101000;
		#400 //-5.2667827e+36 * -2.1853907e-25 = 1150997800000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001101011001111110011000001101;
		b = 32'b10011001101000010111110101001100;
		correct = 32'b10100111100100100100100100101110;
		#400 //243163340.0 * -1.6697617e-23 = -4.060248e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110001001010100100001011110011;
		b = 32'b10000001000010011111100110111011;
		correct = 32'b00110010101101111000011111010111;
		#400 //-8.430942e+29 * -2.53421e-38 = 2.1365777e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001001010110111111100001111010;
		b = 32'b11111100110000110010100101010011;
		correct = 32'b01000110101001111011000111000111;
		#400 //-2.6478e-33 * -8.1066883e+36 = 21464.889
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101001101111111101100010100110;
		b = 32'b00110001001011010000101100101000;
		correct = 32'b01011011100000011010110111000100;
		#400 //2.899099e+25 * 2.5181155e-09 = 7.300266e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101101111000000001010011011101;
		b = 32'b11100011110110111010101011000000;
		correct = 32'b01010010010000000100011101001111;
		#400 //-2.5475117e-11 * -8.1042816e+21 = 206457520000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110011110001110011110010111000;
		b = 32'b00101111100010001000111101001100;
		correct = 32'b00100011110101001000111110010000;
		#400 //9.277704e-08 * 2.4840074e-10 = 2.3045887e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001000010110110011100011010000;
		b = 32'b01001000111011010111111000011100;
		correct = 32'b00010001110010110101111110010111;
		#400 //6.59697e-34 * 486384.88 = 3.2086665e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101000011011011101010100001110;
		b = 32'b00000011001001000101111111101000;
		correct = 32'b00101100000110001011010110010111;
		#400 //4.492524e+24 * 4.8305363e-37 = 2.1701302e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010100101110000000011011110111;
		b = 32'b01000010110000111011010101000001;
		correct = 32'b01011000000011001010111110011010;
		#400 //6323126700000.0 * 97.85401 = 618743300000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101000000000011011110000101011;
		b = 32'b00101111010001111010001110011010;
		correct = 32'b11010111110010100101100001011101;
		#400 //-2.4506255e+24 * 1.8157068e-10 = -444961730000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000101110010010110111010110011;
		b = 32'b01010000010000100111010111001101;
		correct = 32'b10010110100110010000001010010101;
		#400 //-1.8942614e-35 * 13050000000.0 = -2.4720113e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111111010110100110111001101010;
		b = 32'b00000100001001101100110100110011;
		correct = 32'b11000100000011100101001010101111;
		#400 //-2.90345e+38 * 1.9607429e-36 = -569.29193
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110000111011010110000111111100;
		b = 32'b11001011000110000101111111110111;
		correct = 32'b11111100100011010100101100101010;
		#400 //5.8773123e+29 * -9986039.0 = -5.869107e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010100101011001001001111110101;
		b = 32'b00010001110111010101100011000100;
		correct = 32'b10100111000101010011011110010001;
		#400 //-5929733500000.0 * 3.4922358e-28 = -2.0708026e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001000110010011111100011000000;
		b = 32'b10010010000011010010010011001001;
		correct = 32'b10011011010111101011011000001111;
		#400 //413638.0 * -4.4537096e-28 = -1.8422236e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100111010010000111111111001001;
		b = 32'b10011101100010101100000110010110;
		correct = 32'b00000101010110010101100100000000;
		#400 //-2.7824848e-15 * -3.672846e-21 = 1.0219638e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110111101100010000101001000111;
		b = 32'b10000100110110001101011101001101;
		correct = 32'b00111101000101011111010110010001;
		#400 //-7.1816015e+33 * -5.097908e-36 = 0.036611143
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000001011101110101101011001010;
		b = 32'b11100111000010001011001001110101;
		correct = 32'b11101001000001000001010010101001;
		#400 //15.459665 * -6.455338e+23 = -9.979736e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111100100110001011100001101110;
		b = 32'b00101110001111101111101000010001;
		correct = 32'b10101011011000111101110000100000;
		#400 //-0.01864263 * 4.3423102e-11 = -8.0952085e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110110110000101111111111110110;
		b = 32'b00001010111001011011111111000101;
		correct = 32'b11000010001011110000000100001010;
		#400 //-1.9775334e+33 * 2.2124034e-32 = -43.751015
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000010110101011101100010010000;
		b = 32'b11110100010100110100001101111010;
		correct = 32'b00110111101100000111100111011100;
		#400 //-3.1421838e-37 * -6.69521e+31 = 2.103758e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010111001101111100100101101100;
		b = 32'b00110110111010111000000010000100;
		correct = 32'b11001110101010010001001000101010;
		#400 //-202075730000000.0 * 7.018507e-06 = -1418270000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011001010000100010011110001010;
		b = 32'b10110110111001111100100111100001;
		correct = 32'b10010000101011111100101011001001;
		#400 //1.003755e-23 * -6.9078383e-06 = -6.933777e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110001010010001110001111110010;
		b = 32'b10100010010110101010100011010100;
		correct = 32'b10010100001010111001011010011000;
		#400 //2.9233402e-09 * -2.9633886e-18 = -8.662993e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111101110111010000001010101110;
		b = 32'b00001100110011110100011100011001;
		correct = 32'b00001011001100101111001010001100;
		#400 //0.10791527 * 3.193619e-31 = 3.4464025e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010101100111010100001001101001;
		b = 32'b11011101001000101100011010100000;
		correct = 32'b00110011010001111111110000010100;
		#400 //-6.351657e-26 * -7.330774e+17 = 4.6562562e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111011011111100000101111001111;
		b = 32'b10110010010000100111001101000010;
		correct = 32'b01101110010000001111011101010100;
		#400 //-1.3190829e+36 * -1.1318493e-08 = 1.4930031e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110111101010110010101011010111;
		b = 32'b00100111111000010100001110001111;
		correct = 32'b00100000000101101001110111010011;
		#400 //2.0404737e-05 * 6.2523292e-15 = 1.2757714e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001110000111110111110110000011;
		b = 32'b00100100101011000001000000000110;
		correct = 32'b10110011010101100110010010011111;
		#400 //-668950700.0 * 7.4620254e-17 = -4.9917272e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001010110101000100100001110100;
		b = 32'b01001001001111111110111111101011;
		correct = 32'b10010100100111110010100100000001;
		#400 //-2.0442111e-32 * 786174.7 = -1.607107e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110010001110000110111110000010;
		b = 32'b00011101111100000101101000011010;
		correct = 32'b10010000101011010010100101110100;
		#400 //-1.07355635e-08 * 6.3620634e-21 = -6.8300337e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000011111010001010110010100110;
		b = 32'b10100010000000101101101111001001;
		correct = 32'b10100110011011011101111011011101;
		#400 //465.34882 * -1.7734639e-18 = -8.252793e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011100000011001101011011011111;
		b = 32'b00001010011001010011100101101010;
		correct = 32'b10100110111111000011011110010111;
		#400 //-1.58571e+17 * 1.1036747e-32 = -1.750108e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101101100100101001110001010001;
		b = 32'b10011000001111110100110110101110;
		correct = 32'b01000110010110110001111000111010;
		#400 //-5.6717233e+27 * -2.472539e-24 = 14023.557
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110101100001011010110011011000;
		b = 32'b00011001010111001000111010000101;
		correct = 32'b00001111011001100101010111101010;
		#400 //9.959576e-07 * 1.1402515e-23 = 1.1356422e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100111110001110101000001000001;
		b = 32'b00011010111011010110001111010100;
		correct = 32'b10000011001110001101001100000101;
		#400 //-5.5320607e-15 * 9.8182184e-23 = -5.431498e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010000111100111000101011100011;
		b = 32'b11011110010101111101011100110111;
		correct = 32'b01101111110011010101011001100011;
		#400 //-32687725000.0 * -3.88824e+18 = 1.2709772e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011101110101001111010010000011;
		b = 32'b00111000000111001001001000011100;
		correct = 32'b11010110100000100011111010001011;
		#400 //-1.9181292e+18 * 3.7329373e-05 = -71602570000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011101010100100000001100110101;
		b = 32'b10101010010010111010010010110100;
		correct = 32'b10001000001001110000111110101001;
		#400 //2.7794927e-21 * -1.8087165e-13 = -5.0273143e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100011110011001001010111010100;
		b = 32'b11000110101001111100100010000110;
		correct = 32'b01101011000001100001010111111101;
		#400 //-7.547864e+21 * -21476.262 = 1.620999e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001111011001000010000100111101;
		b = 32'b01000101011011101011011001111101;
		correct = 32'b01010101010101001011100110000110;
		#400 //3827383600.0 * 3819.4055 = 14618330000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110100010011010011001100110000;
		b = 32'b11101010010100100001011011010110;
		correct = 32'b01011111001010000110011001001011;
		#400 //-1.9110735e-07 * -6.3495565e+25 = 1.2134469e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011010110011010101001110110001;
		b = 32'b10111001100010011001111101011101;
		correct = 32'b01010100110111001100001100110111;
		#400 //-2.8897195e+16 * -0.0002624941 = 7585343700000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001111101001001001100110101011;
		b = 32'b10110011110111011011010001011001;
		correct = 32'b10000100000011101000110010011110;
		#400 //1.623084e-29 * -1.03239195e-07 = -1.6756588e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100010011011010010000001011000;
		b = 32'b11010001001111000110111100011110;
		correct = 32'b10110100001011101000101010101101;
		#400 //3.2136612e-18 * -50582380000.0 = -1.6255463e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110010100100011110111110011101;
		b = 32'b10010001101111011000001000110010;
		correct = 32'b00000100110110000001000000111110;
		#400 //-1.6989185e-08 * -2.9899181e-28 = 5.0796272e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100110101001001000011101010010;
		b = 32'b11010000100001111110111110111111;
		correct = 32'b01110111101011101011101011100011;
		#400 //-3.8848216e+23 * -18245090000.0 = 7.087892e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100111101111110001111001100101;
		b = 32'b01000101000110000110110101110100;
		correct = 32'b11101101011000111001011110000101;
		#400 //-1.8050654e+24 * 2438.8408 = -4.402267e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100001000110010010110101101111;
		b = 32'b11001001110000000010000001100111;
		correct = 32'b10101011011001011110101011101101;
		#400 //5.1898547e-19 * -1573900.9 = -8.168317e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110100111011100100010000010000;
		b = 32'b00001000010111111011110000010110;
		correct = 32'b00111101110100000011110001011000;
		#400 //1.5101894e+32 * 6.7327715e-34 = 0.1016776
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101111101011111111100100101011;
		b = 32'b10101110101000010010000111100000;
		correct = 32'b10011110110111011000010111111010;
		#400 //3.200936e-10 * -7.32745e-11 = -2.3454697e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000001000011011110001111100011;
		b = 32'b11011011101100011011001001011001;
		correct = 32'b00011101010001001111101011010011;
		#400 //-2.606111e-38 * -1.0003433e+17 = 2.6070057e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000100001111110110110101110110;
		b = 32'b11010011111000100000110000101000;
		correct = 32'b01011000101010010000011110111001;
		#400 //-765.7103 * -1941733100000.0 = 1486805100000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101100100000010110100001011100;
		b = 32'b00011011001010100011111001000000;
		correct = 32'b01001000001011000001110110001001;
		#400 //1.251554e+27 * 1.4082184e-22 = 176246.14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100010000111111100110010101000;
		b = 32'b00001111011101011110001011111011;
		correct = 32'b00110010000110010111110010001100;
		#400 //7.3694484e+20 * 1.21231475e-29 = 8.934091e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000100011100111101101100101101;
		b = 32'b11101000110010101000111110110011;
		correct = 32'b10101101110000001111001111010011;
		#400 //2.8665153e-36 * -7.6525505e+24 = -2.1936153e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000111001000011010111101011101;
		b = 32'b00000100010101100010100111011100;
		correct = 32'b10001100000001110100001100001000;
		#400 //-41391.363 * 2.51748e-36 = -1.0420193e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100111000000111110111110000;
		b = 32'b00111011000010000100010011101000;
		correct = 32'b01000000011011101111111010101001;
		#400 //1795.9355 * 0.0020793024 = 3.7342932
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101011111001101100001000100111;
		b = 32'b00011110110111101001100000111011;
		correct = 32'b10001011010010001010010110010110;
		#400 //-1.6396371e-12 * 2.3568125e-20 = -3.8643172e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001011011000001010110010100001;
		b = 32'b11001111010000010010000111011000;
		correct = 32'b00011011001010010111111111011001;
		#400 //-4.3270702e-32 * -3240220700.0 = 1.4020662e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010001101111010111001000100001;
		b = 32'b01011010011111010111101010101000;
		correct = 32'b11101100101110111001010010001111;
		#400 //-101707950000.0 * 1.7837008e+16 = -1.8141654e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101010101000110101101110101011;
		b = 32'b00000001101101110101110110101000;
		correct = 32'b00101100111010100000010010010101;
		#400 //9.87439e+25 * 6.7357973e-38 = 6.6511887e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111110101100110011000100001010;
		b = 32'b10101000101101100111000000010101;
		correct = 32'b11100111111111110110011010100011;
		#400 //1.1909322e+38 * -2.0254667e-14 = -2.4121935e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100000010100111000000011001000;
		b = 32'b10110000001000011000110101100010;
		correct = 32'b11010001000001010111100011001101;
		#400 //6.0961604e+19 * -5.8772376e-10 = -35828584000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100100010000001110010000000110;
		b = 32'b00110100000010001111110000111100;
		correct = 32'b11011000110011100110111001100010;
		#400 //-1.4232823e+22 * 1.275775e-07 = -1815787900000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111010111110111011101010100010;
		b = 32'b01110100001111000001111011000111;
		correct = 32'b01101111101110001111101101010011;
		#400 //0.0019205401 * 5.961768e+31 = 1.1449815e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101000010001001111010001011111;
		b = 32'b00101110010000110110111010100100;
		correct = 32'b00010111000101100101101101000100;
		#400 //1.0933175e-14 * 4.4436135e-11 = 4.8582807e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111101001010111001001010111010;
		b = 32'b00111100010110000101011011000111;
		correct = 32'b10111010000100001111110111110110;
		#400 //-0.041887976 * 0.013204283 = -0.0005531007
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101101110001010110110111101110;
		b = 32'b10111100000111101000011001111110;
		correct = 32'b11101010011101001000001100100011;
		#400 //7.6376805e+27 * -0.00967562 = -7.3899294e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010010101110101000110111100111;
		b = 32'b01011101100111100000001100110110;
		correct = 32'b00110000111001100100101111010111;
		#400 //1.1773232e-27 * 1.4232505e+18 = 1.6756257e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110110101100101101100101100111;
		b = 32'b01110011110110001101010101010001;
		correct = 32'b01101011000101110111110001110110;
		#400 //5.3301223e-06 * 3.4358603e+31 = 1.8313555e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001001111100011101100100101000;
		b = 32'b10000110011110000001001011010000;
		correct = 32'b10010000111010100101110000100101;
		#400 //1981221.0 * -4.6657437e-35 = -9.24387e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000011110110011110100001100111;
		b = 32'b01110100011111001110010110110100;
		correct = 32'b01111000110101110100010001001011;
		#400 //435.81564 * 8.0146347e+31 = 3.492903e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000001001000101010110101101010;
		b = 32'b11101100000010110101110110100000;
		correct = 32'b10101101101100010001111101001110;
		#400 //2.987912e-38 * -6.739313e+26 = -2.0136472e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011100011110110101000110110101;
		b = 32'b01010011000001001110100100100001;
		correct = 32'b10110000000000100111101011111111;
		#400 //-8.3154537e-22 * 570846940000.0 = -4.746851e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100100100100110111011000001110;
		b = 32'b01110011001010001101110001010100;
		correct = 32'b01011000010000101000100011000110;
		#400 //6.395108e-17 * 1.337852e+31 = 855570800000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110100101110000110110011011100;
		b = 32'b00000100010000000100001011111001;
		correct = 32'b00111001100010101000000111100100;
		#400 //1.1689338e+32 * 2.2600244e-36 = 0.00026418187
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100101110101011011000010010110;
		b = 32'b11101000101111011011111001111111;
		correct = 32'b01001111000111100110001001100010;
		#400 //-3.706927e-16 * -7.1683304e+24 = 2657247700.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100110100110101001001100011111;
		b = 32'b01100111110011110100110010110001;
		correct = 32'b01001110111110100101011010001001;
		#400 //1.0725774e-15 * 1.9578891e+24 = 2099987600.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100111011000100110010011110111;
		b = 32'b01000110110000011001010111011110;
		correct = 32'b11101110101010110011001010100111;
		#400 //-1.0691173e+24 * 24778.934 = -2.6491586e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100010010000101100110011010000;
		b = 32'b10010000001101101000000100010000;
		correct = 32'b10110011000010101101111111010001;
		#400 //8.9835666e+20 * -3.5992597e-29 = -3.233419e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000111100100100101101001001111;
		b = 32'b10100010011000000011011001111001;
		correct = 32'b00101010100000000010111000101001;
		#400 //-74932.62 * -3.0386498e-18 = 2.2769398e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111010100101001001100111101000;
		b = 32'b00111111001010111100000111000011;
		correct = 32'b11111010010001110110011010001110;
		#400 //-3.8579076e+35 * 0.6709253 = -2.5883678e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010010110001011100111010011100;
		b = 32'b11011110101001111001110100111111;
		correct = 32'b11110010000000011000001101001000;
		#400 //424787440000.0 * -6.0389395e+18 = -2.5652656e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010011100010010000011000001000;
		b = 32'b11110000010111010010100100100011;
		correct = 32'b11000100011011001100000001110011;
		#400 //3.458961e-27 * -2.7378367e+29 = -947.007
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011000111010101010101011111111;
		b = 32'b11000011001011101010101111010010;
		correct = 32'b00011100101000000001110110111010;
		#400 //-6.0660244e-24 * -174.67117 = 1.0595596e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101010011111010111001110111110;
		b = 32'b00010110111011011011100101011101;
		correct = 32'b11000001111010110101101110101100;
		#400 //-7.6601202e+25 * 3.8406396e-25 = -29.419762
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111110110101000010000101010000;
		b = 32'b00101010111011111110011001100101;
		correct = 32'b01101010010001101100101000000011;
		#400 //1.4098465e+38 * 4.2614797e-13 = 6.008032e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010010110100011100100110110101;
		b = 32'b11100010101110100000111110110101;
		correct = 32'b00110110000110000111100101101101;
		#400 //-1.3239479e-27 * -1.7161131e+21 = 2.2720444e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011100110111101000110110001000;
		b = 32'b11100011110100011110110011011101;
		correct = 32'b01000001001101100111111101110111;
		#400 //-1.4727313e-21 * -7.7448746e+21 = 11.406119
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010001100011001101110110101111;
		b = 32'b01100000001010001111010111100010;
		correct = 32'b10110010001110011111000110001111;
		#400 //-2.2224728e-28 * 4.8699543e+19 = -1.0823341e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011001000000100000011110011010;
		b = 32'b11101110111001011010111100111100;
		correct = 32'b11001000011010010101001110011101;
		#400 //6.7223776e-24 * -3.5541956e+28 = -238926.45
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011000110100100000010101111011;
		b = 32'b00101110100000110011100110001110;
		correct = 32'b01000111110101110101000000001011;
		#400 //1847367800000000.0 * 5.967414e-11 = 110240.086
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010101101011001101011111001101;
		b = 32'b10101111010010110011001101100100;
		correct = 32'b00000101100010010011000111010010;
		#400 //-6.981072e-26 * -1.8481e-10 = 1.2901719e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100010001110000111000000110001;
		b = 32'b00100011101101000001100110000110;
		correct = 32'b00000110100000011100000101000110;
		#400 //2.4996044e-18 * 1.9526449e-17 = 4.8808397e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001100000110111010000101101110;
		b = 32'b00110110101110000110111010111100;
		correct = 32'b01000011011000000011111010110001;
		#400 //40797624.0 * 5.4965185e-06 = 224.24489
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001011110110000010010010011011;
		b = 32'b01010011100001010000101001101111;
		correct = 32'b10011111111000001010011110100111;
		#400 //-8.325525e-32 * 1142811400000.0 = -9.514505e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000000000110100001000010010101;
		b = 32'b11011000001010111111011001000111;
		correct = 32'b00011000000011000001000100110110;
		#400 //-2.393671e-39 * -756296970000000.0 = 1.8103265e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110010000101100100111101100100;
		b = 32'b10100011101100111110010010100110;
		correct = 32'b00010110010100110011111110000110;
		#400 //-8.7492005e-09 * -1.9504055e-17 = 1.7064489e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111111100111001111010010011101;
		b = 32'b10001101011100000001100110001111;
		correct = 32'b10001101100100110011010011111111;
		#400 //1.226215 * -7.3986475e-31 = -9.072333e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110001011101100100001011101011;
		b = 32'b00011000001000101000100010100101;
		correct = 32'b10001010000111000101100111001011;
		#400 //-3.583575e-09 * 2.1006997e-24 = -7.528015e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101101000100100100111010101100;
		b = 32'b00100010010110011011100011101011;
		correct = 32'b11001111111110001101110010111101;
		#400 //-2.829995e+27 * 2.9506879e-18 = -8350431700.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010010001010110001101100110011;
		b = 32'b01111111010001010010110100001111;
		correct = 32'b01010010000000111100101000001100;
		#400 //5.399161e-28 * 2.6209187e+38 = 141507620000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101001000001000011001110101011;
		b = 32'b11111010101001110001000111100110;
		correct = 32'b11100100001011001000110111100110;
		#400 //2.9354703e-14 * -4.337383e+35 = -1.2732259e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011111001010111100101011100111;
		b = 32'b00000000111000110111101101001111;
		correct = 32'b00100000100110001010011110101010;
		#400 //1.237896e+19 * 2.0890892e-38 = 2.5860752e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110000110011001011100011101011;
		b = 32'b10101101010110011111111111110011;
		correct = 32'b11011110101011100101010101101110;
		#400 //5.0686795e+29 * -1.2391854e-11 = -6.281034e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100101101111100011001100100011;
		b = 32'b01010101000110010011111010010110;
		correct = 32'b01111011011000111011011000011111;
		#400 //1.1227412e+23 * 10530880000000.0 = 1.18234524e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111100100101110010111001010101;
		b = 32'b01100010111101001100001110100101;
		correct = 32'b01100000000100001000101110110011;
		#400 //0.01845471 * 2.2575516e+21 = 4.166246e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010111100100010111101100011;
		b = 32'b10111110111100100001101010110001;
		correct = 32'b00111010011001010000101000001100;
		#400 //-0.0018477257 * -0.4728599 = 0.0008737154
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000010001111000011011100000101;
		b = 32'b11110010110111111010110101010100;
		correct = 32'b10110101101001000111001101011100;
		#400 //1.3827848e-37 * -8.8607613e+30 = -1.2252526e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010100110010101110100001111111;
		b = 32'b10100001100101101011001000100101;
		correct = 32'b00110110111011101110001011011011;
		#400 //-6971872000000.0 * -1.021155e-18 = 7.119362e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100110101010111100000100001001;
		b = 32'b00110010000000001100011001111100;
		correct = 32'b11011001001011001100101101011110;
		#400 //-4.0554277e+23 * 7.495711e-09 = -3039831300000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011100011001100001110010011101;
		b = 32'b11011001110011100011100100000001;
		correct = 32'b10110110101110010101111001000100;
		#400 //7.61376e-22 * -7255815000000000.0 = -5.5244036e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100001110100110001000000000101;
		b = 32'b00110011011010100010000010001101;
		correct = 32'b11010101110000010000011101111011;
		#400 //-4.8667717e+20 * 5.4511975e-08 = -26529734000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011010100010100100001101011111;
		b = 32'b01100000110101110001111100100110;
		correct = 32'b10111011111010000101111011001111;
		#400 //-5.7184306e-23 * 1.240092e+20 = -0.00709138
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010110011111100110011001110011;
		b = 32'b00011001101101101101011001011110;
		correct = 32'b00110000101101011011000111011101;
		#400 //69928992000000.0 * 1.8904941e-23 = 1.3220035e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011101001010011111101010100111;
		b = 32'b10110010010101101101000110000101;
		correct = 32'b01010000000011101010001010100110;
		#400 //-7.6551786e+17 * -1.2504079e-08 = 9572096000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110011000000001101011111111;
		b = 32'b11111000001111101001111001001001;
		correct = 32'b11110111001001101101111010011010;
		#400 //0.21885298 * -1.5464794e+34 = -3.3845163e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000100100010011100010010111100;
		b = 32'b01111010010010101010011101101111;
		correct = 32'b00111111010110100001111010101111;
		#400 //3.2389217e-36 * 2.6305998e+35 = 0.8520307
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101101010001011110100011111011;
		b = 32'b10011101101101111001010111000001;
		correct = 32'b01001011100011011110110101010001;
		#400 //-3.8281377e+27 * -4.859454e-21 = 18602658.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010000001010011011100011100001;
		b = 32'b00000101110011001001010110010000;
		correct = 32'b10010110100001111010001001111011;
		#400 //-11389863000.0 * 1.9239008e-35 = -2.1912966e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110111000011010010010101001;
		b = 32'b10011110010000100011111001101011;
		correct = 32'b00010101101010110011010111001100;
		#400 //-6.7246915e-06 * -1.0283182e-20 = 6.9151226e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110101101000100000010110000100;
		b = 32'b00010011100000011101010101110100;
		correct = 32'b11001001101001000101011110111111;
		#400 //-4.107734e+32 * 3.277466e-27 = -1346295.9
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100011100111110101101111010001;
		b = 32'b00111001000011000011110100010111;
		correct = 32'b01011101001011101001100001111011;
		#400 //5.879297e+21 * 0.00013374198 = 7.863088e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111010001000100110110100110011;
		b = 32'b11011011011000001110101010010001;
		correct = 32'b11010110000011101011010001100000;
		#400 //0.00061960815 * -6.3308303e+16 = -39226340000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001100101110100001010101100000;
		b = 32'b00000100101011111011000111100000;
		correct = 32'b10010001111111110110101111010000;
		#400 //-97561340.0 * 4.1305655e-36 = -4.029835e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011101010111111010101000100000;
		b = 32'b01100100000110110100111101001011;
		correct = 32'b01000010000001111011000101001000;
		#400 //2.9601757e-21 * 1.1459836e+22 = 33.923126
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110010011100101100001010001100;
		b = 32'b11000110110001101100100111011011;
		correct = 32'b10111001101111001000000111100011;
		#400 //1.4130489e-08 * -25444.928 = -0.00035954927
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111010010101000111110000000111;
		b = 32'b11100001001010100111010110001101;
		correct = 32'b11011100000011010111101111101110;
		#400 //0.000810564 * -1.9652606e+20 = -1.5929694e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001010000000011010100101011001;
		b = 32'b01001001111001111111010000110001;
		correct = 32'b11010100011010101111011011111011;
		#400 //-2124374.2 * 1900166.1 = -4036664000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010110011011001000110111111010;
		b = 32'b11001011001011011110111001010110;
		correct = 32'b10100010001000001011100000101101;
		#400 //1.9108728e-25 * -11398742.0 = -2.1781545e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111011001011110011011111011100;
		b = 32'b10101110111001001111011110101011;
		correct = 32'b00101010100111001011011101000100;
		#400 //-0.0026736176 * -1.0412234e-10 = 2.7838333e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101011010010100100000111011110;
		b = 32'b10110100111010101110010110000101;
		correct = 32'b10100000101110011001010110001011;
		#400 //7.1856225e-13 * -4.3752894e-07 = -3.1439178e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011111100111111001000010111100;
		b = 32'b01011001111111001001011110000111;
		correct = 32'b10111010000111010111000011101100;
		#400 //-6.757856e-20 * 8887287500000000.0 = -0.00060059014
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100110110000001111001011101011;
		b = 32'b10011111110011001011110101111000;
		correct = 32'b11000111000110100101000001100001;
		#400 //4.555877e+23 * -8.671081e-20 = -39504.38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000101001010110101011110000110;
		b = 32'b10101010111111101000001011111001;
		correct = 32'b10110000101010100101100010000000;
		#400 //2741.4702 * -4.5210344e-13 = -1.2394281e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001100011101000011000000011010;
		b = 32'b00101010011100100100111100110010;
		correct = 32'b00110111011001110010000100000011;
		#400 //64012390.0 * 2.1521394e-13 = 1.3776359e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111100101111011011000110111100;
		b = 32'b00111101100010100100101000111011;
		correct = 32'b11111010110011001111000110100001;
		#400 //-7.879592e+36 * 0.067524396 = -5.320647e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001001111100011000111100111110;
		b = 32'b11010101000011100001010111100001;
		correct = 32'b01011111100001100001001000011001;
		#400 //-1978855.8 * -9764039000000.0 = 1.9321623e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000110000011101010010111001010;
		b = 32'b10100100101010001111110100000100;
		correct = 32'b00101011001111000101001110010001;
		#400 //-9129.447 * -7.328701e-17 = 6.690699e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010010111111001101110001110100;
		b = 32'b11010100110110011000100010100000;
		correct = 32'b00101000010101101101110111010001;
		#400 //-1.5957782e-27 * -7474400700000.0 = 1.1927485e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110010000100100001100101100011;
		b = 32'b00100000110010011101001110110111;
		correct = 32'b00010011011001100101110110000100;
		#400 //8.504091e-09 * 3.4190826e-19 = 2.9076188e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010001111010110100101011011101;
		b = 32'b01010100101000100010000111010011;
		correct = 32'b11100111000101010000010001110110;
		#400 //-126321660000.0 * 5570817400000.0 = -7.037149e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111001001111111000111110001111;
		b = 32'b00000010111001100100001100010101;
		correct = 32'b00111100101011000100110100101101;
		#400 //6.2165026e+34 * 3.3833966e-37 = 0.021032894
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101110110001010000001000110010;
		b = 32'b01101010000011011101001111100000;
		correct = 32'b01011001010110100100101010000101;
		#400 //8.958913e-11 * 4.2864773e+25 = 3840217500000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100101111000001110100110101001;
		b = 32'b01101111010111100101010011001100;
		correct = 32'b11010101110000110101010100100000;
		#400 //-3.901614e-16 * 6.8808185e+28 = -26846297000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000001011111110010011100010011;
		b = 32'b11001110100011110000001000100000;
		correct = 32'b11010000100011101000100011110010;
		#400 //15.94704 * -1199640600.0 = -19130716000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110010011000000100011011110110;
		b = 32'b01100101001101001011101111001100;
		correct = 32'b11011000000111100101011001101100;
		#400 //-1.3054651e-08 * 5.334314e+22 = -696376070000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110110111001010011101000110111;
		b = 32'b10111010111011001001111011100010;
		correct = 32'b01110010010100111101111111101111;
		#400 //-2.324642e+33 * -0.0018052722 = 4.1966116e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101110010010000110100011011101;
		b = 32'b10111001110010100010011111010101;
		correct = 32'b10101000100111100100000111101101;
		#400 //4.5567872e-11 * -0.0003855812 = -1.7570115e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100000011001101101011001111010;
		b = 32'b01010100100110011111001101101110;
		correct = 32'b11110101100010101101000110110000;
		#400 //-6.6534466e+19 * 5289712500000.0 = -3.519482e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111100111010111011001100111001;
		b = 32'b01100001011110100010010000011100;
		correct = 32'b01011110111001100100111001000101;
		#400 //0.028771983 * 2.88393e+20 = 8.297639e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000000110000110110110001110011;
		b = 32'b00000101110011001011010001000100;
		correct = 32'b10000111000111000100010000001000;
		#400 //-6.1069884 * 1.9250287e-35 = -1.1756128e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010010000100100011110101011011;
		b = 32'b11001100110010001110110010101111;
		correct = 32'b00011111011001011000111001000111;
		#400 //-4.6145103e-28 * -105342330.0 = 4.8610325e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111110111110100011111011111000;
		b = 32'b00000101000100000011000101001000;
		correct = 32'b11000100100011001111001110011000;
		#400 //-1.6631698e+38 * 6.779899e-36 = -1127.6123
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100010010110010100000110010011;
		b = 32'b01000011011101110111100110111000;
		correct = 32'b10100110010100100000010110010001;
		#400 //-2.9443699e-18 * 247.47546 = -7.286593e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110001100011010101110111110001;
		b = 32'b00010000100000111101100100100001;
		correct = 32'b10000010100100011001110111110010;
		#400 //-4.11432e-09 * 5.200493e-29 = -2.1396491e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101101011011100100001011011110;
		b = 32'b01111011000001011010011111001110;
		correct = 32'b11101000111110001100100111010101;
		#400 //-1.3543581e-11 * 6.93979e+35 = -9.39896e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001110111011011100000101011100;
		b = 32'b11101010111110001000111100101110;
		correct = 32'b11111010011001101101100001001011;
		#400 //1994436100.0 * -1.50244875e+26 = -2.996538e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011010100111101011110011101011;
		b = 32'b11110100011001000011000110111010;
		correct = 32'b01001111100011010111111100010111;
		#400 //-6.565248e-23 * -7.2317643e+31 = 4747833000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011100101101100110000111000000;
		b = 32'b01011000001011100001111001000110;
		correct = 32'b01110101011110000001100000000100;
		#400 //4.106874e+17 * 765780200000000.0 = 3.1449627e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000010100101111101011110110101;
		b = 32'b01011001101000000010110011001011;
		correct = 32'b11011100101111100000001011000101;
		#400 //-75.9213 * 5635656000000000.0 = -4.2786633e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101010011000100101010011100110;
		b = 32'b10100001010001010000010000001100;
		correct = 32'b01001100001011100010111011101001;
		#400 //-6.840454e+25 * -6.675155e-19 = 45661092.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111100100110100101001100000001;
		b = 32'b00000110010000011001110100001011;
		correct = 32'b10000011011010010110111001111111;
		#400 //-0.018838407 * 3.6414643e-35 = -6.859939e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100110011101110010010101011001;
		b = 32'b11000010100001111100101010110000;
		correct = 32'b10101001100000110001100001011111;
		#400 //8.5745955e-16 * -67.895874 = -5.8217964e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101000101011100011111001010010;
		b = 32'b00100011010110100000001100111001;
		correct = 32'b01001100100101000110001101000011;
		#400 //6.582731e+24 * 1.1818486e-17 = 77797910.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110111101000010111001111000000;
		b = 32'b11000100100100001101001010100001;
		correct = 32'b11111100101101101010101111100101;
		#400 //6.549277e+33 * -1158.5822 = -7.587876e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100011101110100000101001000110;
		b = 32'b10101001000000101101100100110110;
		correct = 32'b01001101001111100010111000100011;
		#400 //-6.8636694e+21 * -2.90542e-14 = 199418420.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101011011011011101001111110101;
		b = 32'b11000100000110010111011100111111;
		correct = 32'b01110000000011101001001001110101;
		#400 //-2.8751636e+26 * -613.8632 = 1.764957e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001011001111001001111101101010;
		b = 32'b10111000101100000110111001101010;
		correct = 32'b11000100100000011111111011110011;
		#400 //12361578.0 * -8.4129e-05 = -1039.9672
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111111111110110110011011111111;
		b = 32'b10010100001011100110101100111111;
		correct = 32'b11111111111110110110011011111111;
		#400 //nan * -8.8059056e-27 = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100101000100111110001110000011;
		b = 32'b11011011101100110111100010100010;
		correct = 32'b01000001010011110101101110001010;
		#400 //-1.2827302e-16 * -1.0103332e+17 = 12.959848
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011010000001110011111111101000;
		b = 32'b01010110001100011111011110101010;
		correct = 32'b00110000101111000000110000010000;
		#400 //2.796897e-23 * 48919317000000.0 = 1.3682229e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000000100001101000010100110011;
		b = 32'b00000001101100101111110010011011;
		correct = 32'b10000010101111000001101010110100;
		#400 //-4.2037597 * 6.5749344e-38 = -2.7639444e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011111101111111110010110100010;
		b = 32'b11101110100111111011001110111011;
		correct = 32'b11001110111011110110110010110011;
		#400 //8.127154e-20 * -2.4712699e+28 = -2008439200.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110011110101001000010000001110;
		b = 32'b11110111101001111111111010000101;
		correct = 32'b01101100000010110111010101101111;
		#400 //-9.89604e-08 * -6.814655e+33 = 6.74381e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111101001010010000111100110110;
		b = 32'b10101111010111110111010001110100;
		correct = 32'b01101101000100111001000100101000;
		#400 //-1.4044907e+37 * -2.0323104e-10 = 2.8543612e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011111001001011101110000100001;
		b = 32'b00000111100111011011101100111111;
		correct = 32'b00100111010011000110001010100010;
		#400 //1.1951464e+19 * 2.3732788e-34 = 2.8364156e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100110110111100010110111010100;
		b = 32'b10111111010011100100000001011001;
		correct = 32'b01100110101100110000000010111001;
		#400 //-5.2460537e+23 * -0.80566937 = 4.2265847e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010011001001000000110110101110;
		b = 32'b11110000110111011111010110100010;
		correct = 32'b01000100100011100011110100111000;
		#400 //-2.0706455e-27 * -5.495451e+29 = 1137.9131
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011101010100001011011100100010;
		b = 32'b00110010110100010101101001001111;
		correct = 32'b00010000101010101010111100100100;
		#400 //2.7623248e-21 * 2.437187e-08 = 6.7323024e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111000111001010111110111110110;
		b = 32'b10101000101010000100011011000101;
		correct = 32'b01100010000101101101101000011010;
		#400 //-3.7237212e+34 * -1.8682438e-14 = 6.956819e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001000010101100001111100010001;
		b = 32'b11101001100011100101000101001101;
		correct = 32'b10110010011011100001001001110111;
		#400 //6.44348e-34 * -2.1506425e+25 = -1.3857622e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110110101100101010101001100011;
		b = 32'b10001100100000100111111100001101;
		correct = 32'b10000011101101100010011001100100;
		#400 //5.324649e-06 * -2.0106137e-31 = -1.0705813e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010101101000111001010110000111;
		b = 32'b00010110010000000011110110010010;
		correct = 32'b00101100011101011010111011111010;
		#400 //22482826000000.0 * 1.5529065e-25 = 3.4913726e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000001001011001110101100011011;
		b = 32'b11110111000010011100000111000101;
		correct = 32'b11111000101110100001100101101000;
		#400 //10.807399 * -2.794042e+33 = -3.0196329e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101001111000001110101100001110;
		b = 32'b11010011011001110101100010000011;
		correct = 32'b10111101110010110100000111011110;
		#400 //9.988374e-14 * -993622400000.0 = -0.099246725
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101010100000000111011011011000;
		b = 32'b11010000011001011111011010110000;
		correct = 32'b00111011011001101100110000110011;
		#400 //-2.2819832e-13 * -15432598000.0 = 0.0035216927
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111100010010011001101111101100;
		b = 32'b01100011000000000010111010001111;
		correct = 32'b11011111110010011110010101000001;
		#400 //-0.012305241 * 2.3645381e+21 = -2.9096211e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000110101100100011010100110001;
		b = 32'b10111000100101000100100010110100;
		correct = 32'b10111111110011100111001010111001;
		#400 //22810.596 * -7.070732e-05 = -1.612876
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001010010110110010010111110101;
		b = 32'b00011100101100110000101100010010;
		correct = 32'b00100111100110010100010100000100;
		#400 //3590525.2 * 1.1848088e-21 = 4.2540858e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001111010010110111001010101001;
		b = 32'b00101110111101000100000101101010;
		correct = 32'b00111110110000100001110101000101;
		#400 //3413289200.0 * 1.1107455e-10 = 0.37912956
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110101100101100000011110010100;
		b = 32'b10111110101101111010100111010001;
		correct = 32'b11110100110101110100010111100001;
		#400 //3.8037023e+32 * -0.35871747 = -1.3644545e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011011110011100011011100011111;
		b = 32'b11001010101100000000001101000111;
		correct = 32'b10100111000011011100100010001001;
		#400 //3.4115462e-22 * -5767587.5 = -1.9676391e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010001110101010111101000001110;
		b = 32'b00000111101100001010100110001001;
		correct = 32'b00011010000100110101000101001001;
		#400 //114609470000.0 * 2.658118e-34 = 3.046455e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101001011001110100100001100100;
		b = 32'b01011001110011111110101000001111;
		correct = 32'b01000011101110111101011011111111;
		#400 //5.1355093e-14 * 7315334000000000.0 = 375.67966
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001001000110010100101000001111;
		b = 32'b10111110110001110111111000011110;
		correct = 32'b10001000011011101110100000101100;
		#400 //1.8451527e-33 * -0.38963407 = -7.1893437e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101000111010001111111111001000;
		b = 32'b01100100000110000101010010100111;
		correct = 32'b11001101100010101010010011101011;
		#400 //-2.5868102e-14 * 1.124002e+22 = -290757980.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000010010010010111011000000010;
		b = 32'b01011000111100010111111110011100;
		correct = 32'b01011011101111100000110010000100;
		#400 //50.365242 * 2124243000000000.0 = 1.0698801e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100101001010100101011010101110;
		b = 32'b01010101100001010001001110011101;
		correct = 32'b01111011001100010001100000101011;
		#400 //5.027508e+22 * 18289910000000.0 = 9.195267e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011011111011000110100100011110;
		b = 32'b10101100010101100010101000101100;
		correct = 32'b00001000110001011100011011010001;
		#400 //-3.9110855e-22 * -3.043464e-12 = 1.1903248e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100000010101011011011100000011;
		b = 32'b01010010110111110010101100000010;
		correct = 32'b11110011101110100100111001010011;
		#400 //-6.1599123e+19 * 479249630000.0 = -2.9521357e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011001100110000100100101101110;
		b = 32'b01000011011011101111110000010101;
		correct = 32'b10011101100011100010101000111001;
		#400 //-1.574609e-23 * 238.9847 = -3.7630744e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011101011000010100011110010110;
		b = 32'b10101101100110011111000110101111;
		correct = 32'b01001011100001110111100001110111;
		#400 //-1.0145693e+18 * -1.7501415e-11 = 17756398.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001101011000000000100100011001;
		b = 32'b11101000010101001111011111011111;
		correct = 32'b00110110001110100110000001110101;
		#400 //-6.903628e-31 * -4.0228564e+24 = 2.7772305e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001010101000111100001001110011;
		b = 32'b01110000011000011000100111100111;
		correct = 32'b11111011100100000100011000011110;
		#400 //-5366073.5 * 2.7920336e+29 = -1.4982258e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110101001101100101110010000101;
		b = 32'b00110001111111110101000110110010;
		correct = 32'b01100111101101011110000001011011;
		#400 //2.3117054e+32 * 7.4307644e-09 = 1.7177739e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100000111001001010100011001111;
		b = 32'b10000111011100010110001010110100;
		correct = 32'b00101000110101111001101100010100;
		#400 //-1.31813175e+20 * -1.8159831e-34 = 2.393705e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101010111101100011011101001100;
		b = 32'b01101001101100001101011100111000;
		correct = 32'b11010101001010100001010100000011;
		#400 //-4.3736748e-13 * 2.672341e+25 = -11687951000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111011111000010010010110010010;
		b = 32'b10100111001110001111110000101001;
		correct = 32'b11100011101000101011000011000110;
		#400 //2.3380576e+36 * -2.5671826e-15 = -6.002221e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010001011100100010111110100101;
		b = 32'b10100001100111110100011101110110;
		correct = 32'b00110011100101101010111100110010;
		#400 //-65011340000.0 * -1.0793175e-18 = 7.016787e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101011110101010101100010101011;
		b = 32'b11011101010010110100011011011010;
		correct = 32'b11001001101010010110100001011100;
		#400 //1.5159171e-12 * -9.1547716e+17 = -1387787.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111011000001100100111100101110;
		b = 32'b10001001101000111110011110010111;
		correct = 32'b01000101001010111111101111010110;
		#400 //-6.973737e+35 * -3.945861e-33 = 2751.7397
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010000011010000101100101010101;
		b = 32'b01001111110100100000100001101111;
		correct = 32'b11100000101111101010000011101111;
		#400 //-15592674000.0 * 7047536000.0 = -1.0988993e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100010001010011011100001100110;
		b = 32'b11111100010011001110110101010010;
		correct = 32'b01011111000001111101110001000111;
		#400 //-2.300139e-18 * -4.256168e+36 = 9.789778e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001111110101000000010111010010;
		b = 32'b00101111111000001110010100101111;
		correct = 32'b01000000001110100100001011101000;
		#400 //7114302500.0 * 4.0908207e-10 = 2.9103336
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101101011110011101000111100010;
		b = 32'b11011110011100111001011011001110;
		correct = 32'b11001100011011011011010101100100;
		#400 //1.4200615e-11 * -4.3881108e+18 = -62313870.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010100010001101010001001101001;
		b = 32'b00111110101110001001100000101101;
		correct = 32'b11010011100011110011101011001111;
		#400 //-3412513300000.0 * 0.360536 = -1230334000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110010001010011010111000000101;
		b = 32'b11000100011101111110111101001001;
		correct = 32'b10110111001001000101010110000001;
		#400 //9.876662e-09 * -991.73883 = -9.79507e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100011110100000011110010001100;
		b = 32'b10010010011110001011110011001000;
		correct = 32'b00110110110010100101010000110111;
		#400 //-7.682571e+21 * -7.8487693e-28 = 6.029873e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011111010111011000010101000;
		b = 32'b01011110000000010000110111011001;
		correct = 32'b11101010011011011010000110001001;
		#400 //-30892368.0 * 2.3248318e+18 = -7.181956e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010110110001001011011111100110;
		b = 32'b11001001101110101100100000000111;
		correct = 32'b11100001000011111000011101010010;
		#400 //108147060000000.0 * -1530112.9 = -1.654772e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011000100001110101111001101100;
		b = 32'b11110011101101011101001101100001;
		correct = 32'b11001100110000000100101100010001;
		#400 //3.4992024e-24 * -2.8811432e+31 = -100817030.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001101001000010101011100110101;
		b = 32'b11001111111000001111000001100100;
		correct = 32'b00011101100011011100001111001111;
		#400 //-4.9716927e-31 * -7547701000.0 = 3.752485e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100001101111100101111110001100;
		b = 32'b01010011100011011001100000100101;
		correct = 32'b11110101110100101001011110001001;
		#400 //-4.3897078e+20 * 1216285900000.0 = -5.33914e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101011101100000000111001000101;
		b = 32'b10111001110001111001011110100001;
		correct = 32'b11100110000010010100001101011111;
		#400 //4.2567666e+26 * -0.0003806921 = -1.6205175e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001101001100100111100111010101;
		b = 32'b00100100010100011111100001110001;
		correct = 32'b00110010000100100110001010101100;
		#400 //187145550.0 * 4.553009e-17 = 8.520754e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001110111001000000101011100010;
		b = 32'b00001111011100110011100000001111;
		correct = 32'b00011110110110001010100001000100;
		#400 //1912959200.0 * 1.19916215e-29 = 2.2939483e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111111110101001111101111010111;
		b = 32'b10010110111000000010111001110011;
		correct = 32'b10010111001110101000001100000001;
		#400 //1.6639355 * -3.6218465e-25 = -6.026519e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001010111011100011100111000100;
		b = 32'b10100111111001000111111100101100;
		correct = 32'b00110011010101001010000111001010;
		#400 //-7806178.0 * -6.3420592e-15 = 4.9507243e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100110000011010000010111011010;
		b = 32'b01000111101000110100101000101001;
		correct = 32'b11101110001100111110011100101000;
		#400 //-1.664904e+23 * 83604.32 = -1.3919317e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101001001111111111001110110101;
		b = 32'b10111011011001011011111101011110;
		correct = 32'b00100101001011000100010001111110;
		#400 //-4.2621902e-14 * -0.003505669 = 1.4941828e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101110111010011011110110101000;
		b = 32'b10001001010001101100111111101101;
		correct = 32'b00111000101101011000011010001001;
		#400 //-3.6169644e+28 * -2.393115e-33 = 8.655812e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000011100000000001100010001100;
		b = 32'b00100100100001110000100000010010;
		correct = 32'b00101000100001110010000111110111;
		#400 //256.19177 * 5.856059e-17 = 1.500274e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110011010111001100111110110100;
		b = 32'b11110011010011001110111100011101;
		correct = 32'b01100111001100001100001111000010;
		#400 //-5.1411646e-08 * -1.6236547e+31 = 8.347476e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111111011011100101010110011010;
		b = 32'b01011110100000001010011111001011;
		correct = 32'b01011110011011111000111000001000;
		#400 //0.9309937 * 4.635301e+18 = 4.3154358e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000101010011001010010011010001;
		b = 32'b11100010111101001111000010110110;
		correct = 32'b00101000110000111100110110000011;
		#400 //-9.622306e-36 * -2.2591753e+21 = 2.1738475e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100100111010111100011110011011;
		b = 32'b10110111110101011000100100000011;
		correct = 32'b10011101010001001010101101000101;
		#400 //1.0225315e-16 * -2.545538e-05 = -2.6028928e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111111110111100001000100111001;
		b = 32'b01101100001100111100110010100010;
		correct = 32'b11101100100110111111011110001101;
		#400 //-1.7349006 * 8.694563e+26 = -1.5084202e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001011000011010100011011011000;
		b = 32'b01010011101101010001110001100000;
		correct = 32'b10011111010001111110010101111111;
		#400 //-2.720891e-32 * 1555730300000.0 = -4.2329724e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101001101001001011111000100010;
		b = 32'b00010100001010100111100100010011;
		correct = 32'b10111110010110110110100001011001;
		#400 //-2.4895214e+25 * 8.606684e-27 = -0.21426524
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100010011010010111000111001100;
		b = 32'b01011000011011001111110111111010;
		correct = 32'b01111011010110000001110010000001;
		#400 //1.0765728e+21 * 1042302260000000.0 = 1.12211425e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010011010101110110011000100000;
		b = 32'b11101111010000100100110011011110;
		correct = 32'b11000011001000110111110000010001;
		#400 //2.7187167e-27 * -6.013302e+28 = -163.48463
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100101001001100010000010110101;
		b = 32'b01111000110100000000100000000000;
		correct = 32'b01011110100001101111111111000100;
		#400 //1.4409286e-16 * 3.3755e+34 = 4.8638546e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010110111110010000000100100101;
		b = 32'b10010101101100010001110110000000;
		correct = 32'b10101101001011000100011001111100;
		#400 //136891656000000.0 * -7.1536273e-26 = -9.792719e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010110110100001001100111001;
		b = 32'b11110011111010011110100010111001;
		correct = 32'b01101111010001110100000110111110;
		#400 //-0.0016637809 * -3.7064372e+31 = 6.1666994e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110010010110010110110010111;
		b = 32'b10011101001101100111001000100011;
		correct = 32'b10011100000100001100110011111111;
		#400 //0.1984161 * -2.4146507e-21 = -4.7910555e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010100001011011010010110000000;
		b = 32'b11100101110001010101100111100001;
		correct = 32'b11111010100001011101110101010011;
		#400 //2983224000000.0 * -1.1649552e+23 = -3.4753224e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010101101000001010010101001011;
		b = 32'b11011001001011110000111111100000;
		correct = 32'b00101111010110111011010111101001;
		#400 //-6.488427e-26 * -3079723500000000.0 = 1.9982561e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110101000010001000100100010111;
		b = 32'b11110110110010100101001010110110;
		correct = 32'b01101100010101111101000010010010;
		#400 //-5.086344e-07 * -2.0517999e+33 = 1.043616e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010110011100001001110100011011;
		b = 32'b00001010100000001111011100011000;
		correct = 32'b10100001011100100110110110010111;
		#400 //-66139390000000.0 * 1.2418898e-32 = -8.213783e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100001000100101111111010011010;
		b = 32'b11000001001101001111100000110110;
		correct = 32'b10100010110011111101001100010100;
		#400 //4.9803686e-19 * -11.310598 = -5.633095e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010101110010101110101011100000;
		b = 32'b10011010011000010001011101001010;
		correct = 32'b10110000101100100110101011100101;
		#400 //27888766000000.0 * -4.6547722e-23 = -1.2981586e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101111101111111110011001101100;
		b = 32'b11101101000111100001111010100011;
		correct = 32'b11011101011011010000111001011100;
		#400 //3.4906422e-10 * -3.0584793e+27 = -1.0676057e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000001001100010010010011011010;
		b = 32'b11011010100100111011110001101011;
		correct = 32'b01011100010011000111010100010101;
		#400 //-11.071497 * -2.0791995e+16 = 2.3019851e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001110101000010111001100010111;
		b = 32'b01001101001110111011101011101100;
		correct = 32'b11011100011011001100100111101001;
		#400 //-1354337200.0 * 196849340.0 = -2.6660039e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101010100101001001000111001100;
		b = 32'b10111010011001101100011011010101;
		correct = 32'b10100101100001011110111001100010;
		#400 //2.6391248e-13 * -0.0008803432 = -2.3233357e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110001000010111010101111010101;
		b = 32'b11010111000010111011100011101010;
		correct = 32'b11001000100110000111011001100000;
		#400 //2.0324837e-09 * -153626320000000.0 = -312243.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111100001111000100001110001001;
		b = 32'b01010110011101001101000110101100;
		correct = 32'b11010011001101000000101010010000;
		#400 //-0.011490711 * 67295343000000.0 = -773271300000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001010110000000001011101110100;
		b = 32'b01001011110011011101011011010110;
		correct = 32'b10010111000110100111001111111100;
		#400 //-1.849775e-32 * 26979756.0 = -4.9906477e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110001010000100010110110111011;
		b = 32'b11100100011001101111111001101111;
		correct = 32'b11010110001011110011011000010100;
		#400 //2.825671e-09 * -1.704434e+22 = -48161700000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111000010011100010011001100100;
		b = 32'b11100101011000001011000010110100;
		correct = 32'b11011110001101001110111111100011;
		#400 //4.914998e-05 * -6.6316856e+22 = -3.2594723e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001110100000010000011101100111;
		b = 32'b10101010001111001000000101011101;
		correct = 32'b10111001001111100000010101000110;
		#400 //1082373000.0 * -1.6742636e-13 = -0.00018121777
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110001100101001000001010011000;
		b = 32'b10111000000011010011101110010001;
		correct = 32'b11101010001000111101110011111000;
		#400 //1.4707731e+30 * -3.3672495e-05 = -4.95246e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100110100111010100010011011001;
		b = 32'b01011011100000000010011110001011;
		correct = 32'b11000010100111010111010101101111;
		#400 //-1.0912725e-15 * 7.214455e+16 = -78.72936
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011011011010111110100101001000;
		b = 32'b11111011100000000010001111111111;
		correct = 32'b01010111011011000010101110100000;
		#400 //-1.9514122e-22 * -1.3306882e+36 = 259672110000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111111110110101010110011101011;
		b = 32'b10101010011110011011010110100011;
		correct = 32'b01111111110110101010110011101011;
		#400 //nan * -2.217866e-13 = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100101001011111011100111011110;
		b = 32'b11001100011111101010000000001111;
		correct = 32'b00110010001011101100100001001001;
		#400 //-1.5241805e-16 * -66748476.0 = 1.0173673e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100001001101111010001010010000;
		b = 32'b01011101011111110000010000101110;
		correct = 32'b00111111001101101110110111101101;
		#400 //6.221796e-19 * 1.14849143e+18 = 0.71456796
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100110111010011000000001011101;
		b = 32'b10010010001001001111001100110000;
		correct = 32'b00111001100101100111010000001100;
		#400 //-5.5133964e+23 * -5.2049027e-28 = 0.0002869669
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001110001101010111111100000100;
		b = 32'b10010111111110010100000101011100;
		correct = 32'b00100110101100001011011011100001;
		#400 //-761250050.0 * -1.6107747e-24 = 1.2262023e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110001000011111110011100000101;
		b = 32'b11001000011001010011110100010011;
		correct = 32'b11111010000000001101101111111100;
		#400 //7.125703e+29 * -234740.3 = -1.6726895e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011100101111000011110000001100;
		b = 32'b11000101010110000111010101111110;
		correct = 32'b11100010100111110010100100001110;
		#400 //4.2386654e+17 * -3463.3433 = -1.4679953e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101001111101100101001110010101;
		b = 32'b10001000010010110100000101111010;
		correct = 32'b00110010110000111001001101001000;
		#400 //-3.7223807e+25 * -6.116506e-34 = 2.2767964e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110001000011101000001001011;
		b = 32'b00011001001100101011011010001011;
		correct = 32'b10001111111000011110110001101100;
		#400 //-2.4112112e-06 * 9.2392486e-24 = -2.227778e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111010010100111101011110101110;
		b = 32'b10000110011100100101001110011100;
		correct = 32'b01000001010010001000011100010011;
		#400 //-2.7498729e+35 * -4.5576568e-35 = 12.532977
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011000110010001110010010011010;
		b = 32'b00111001010111100111011000011010;
		correct = 32'b10010010101011101001001011101011;
		#400 //-5.1929617e-24 * 0.00021215566 = -1.1017162e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011101000000010011010110101111;
		b = 32'b01001111100001001101010110110000;
		correct = 32'b00101101000001100001011100010001;
		#400 //1.7100762e-21 * 4457193500.0 = 7.62214e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000011010101010101010101110100;
		b = 32'b11001001001001100001101010011101;
		correct = 32'b01001101000010100110101110010111;
		#400 //-213.3338 * -680361.8 = 145144180.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001110100010100110000011000010;
		b = 32'b00111111111100100011010100101101;
		correct = 32'b11001111000000101110110000110110;
		#400 //-1160798500.0 * 1.8922478 = -2196518400.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101101101101000110101011000100;
		b = 32'b00001011110010001111111010100110;
		correct = 32'b10111010000011011010011011100000;
		#400 //-6.9795467e+27 * 7.742035e-32 = -0.00054035895
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000100001100100100110000110011;
		b = 32'b00100000110001111010110011001110;
		correct = 32'b10100101100010110001000110010110;
		#400 //-713.1906 * 3.3826264e-19 = -2.4124573e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101110100001010111000100100110;
		b = 32'b11111011101010011110011111111010;
		correct = 32'b01101010101100010010000100111011;
		#400 //-6.068239e-11 * -1.7644064e+36 = 1.070684e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011000000010011000100010110001;
		b = 32'b11101100010111000101001011111110;
		correct = 32'b11000100111011001011110000011101;
		#400 //1.7775847e-24 * -1.0654224e+27 = -1893.8785
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101101000100111100110110101101;
		b = 32'b00011111010110011111100000101111;
		correct = 32'b10001100111110111011000101000100;
		#400 //-8.401652e-12 * 4.615683e-20 = -3.877936e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100110011010100101001111101010;
		b = 32'b00000011100101011101011111101001;
		correct = 32'b00101010100010010010100001111001;
		#400 //2.7664542e+23 * 8.8070035e-37 = 2.4364172e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110000110111110100110011000000;
		b = 32'b11011110011000100110100011001011;
		correct = 32'b11001111110001010111110100101010;
		#400 //1.6247199e-09 * -4.0786282e+18 = -6626628600.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011001001011001111000001001001;
		b = 32'b11000010111101011011101010111110;
		correct = 32'b10011100101001100000000000011101;
		#400 //8.940717e-24 * -122.86473 = -1.0984988e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110001000101001001101110110001;
		b = 32'b11101001100000010101101110100111;
		correct = 32'b01011011000101100010111101010001;
		#400 //-2.1625335e-09 * -1.954803e+25 = 4.227327e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010010011000111001101101101110;
		b = 32'b11100110100101101001000100000111;
		correct = 32'b00111001100001011101111000000100;
		#400 //-7.182015e-28 * -3.5551513e+23 = 0.0002553315
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001000001000101010000011011111;
		b = 32'b10011011011101010010010001010111;
		correct = 32'b00100100000110111011101100001011;
		#400 //-166531.48 * -2.0277667e-22 = 3.37687e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010001101010011011101000100011;
		b = 32'b11101110011011010011110001000101;
		correct = 32'b11000000100111010100100101001000;
		#400 //2.6778214e-28 * -1.8355202e+28 = -4.9151955
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010011100001001010111000011100;
		b = 32'b10111110101101001111000001111001;
		correct = 32'b01010010101110111000111000011011;
		#400 //-1139713500000.0 * -0.35339716 = 402771500000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110110010111111101010010110101;
		b = 32'b00110101010110001001111101110100;
		correct = 32'b11101100001111010110011011100011;
		#400 //-1.1349574e+33 * 8.0698305e-07 = -9.158914e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011011001011110001110001011111;
		b = 32'b10101010011110100010010101110110;
		correct = 32'b01000110001010110001101101010101;
		#400 //-4.9289315e+16 * -2.2217457e-13 = 10950.833
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011110110010100111001000011110;
		b = 32'b00111000010101010000100010010111;
		correct = 32'b00010111101010000111011110111110;
		#400 //2.143478e-20 * 5.0791157e-05 = 1.0886973e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010111100101110010000101000111;
		b = 32'b01001000101000000011100100010111;
		correct = 32'b10100000101111010010110100000001;
		#400 //-9.766547e-25 * 328136.72 = -3.2047626e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101011011010010111110001101110;
		b = 32'b10010111100111101010010001110100;
		correct = 32'b10000011100100001011000011001001;
		#400 //8.295091e-13 * -1.0252024e-24 = -8.504147e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101000001011110010001111000101;
		b = 32'b11101000110001011000001000100011;
		correct = 32'b11010001100001110001111110001111;
		#400 //9.722208e-15 * -7.4616544e+24 = -72543760000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100001110111111010101011101101;
		b = 32'b01011011111111100111111011100100;
		correct = 32'b01111110010111100101101001110100;
		#400 //5.1574255e+20 * 1.4326832e+17 = 7.388957e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000111100111011100111000100111;
		b = 32'b11101101101111101011000111111000;
		correct = 32'b00110101111010110001100101101011;
		#400 //-2.37439e-34 * -7.377163e+27 = 1.7516262e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111111111010101100011000111110;
		b = 32'b11001101001001111000010011001110;
		correct = 32'b01111111111010101100011000111110;
		#400 //nan * -175656160.0 = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010000100010001100000010011101;
		b = 32'b11100011101000000010111110101111;
		correct = 32'b01110100101010110010001110110110;
		#400 //-18354596000.0 * -5.90983e+21 = 1.0847254e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010100001001011011001011011110;
		b = 32'b11110000100001110001001101010010;
		correct = 32'b01000101001011101101101110101001;
		#400 //-8.3656465e-27 * -3.3443067e+29 = 2797.7288
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110001000010011010000100001011;
		b = 32'b00110011101011001000010011111110;
		correct = 32'b00100101001110010111111101100110;
		#400 //2.0027666e-09 * 8.033565e-08 = 1.6089356e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100000101110001000011011011010;
		b = 32'b00000101100101011100110110010101;
		correct = 32'b10100110110101111111010101011001;
		#400 //-1.0637244e+20 * 1.4087412e-35 = -1.4985124e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001000100110011100001010011100;
		b = 32'b10011101101100001110101110010010;
		correct = 32'b10100110110101001000011010010001;
		#400 //314900.88 * -4.6830386e-21 = -1.4746929e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111111111011011110001000011100;
		b = 32'b01110001101101100001000001001000;
		correct = 32'b01111111111011011110001000011100;
		#400 //nan * 1.8030705e+30 = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101010001111001001111010110101;
		b = 32'b10010101100111001001000111101110;
		correct = 32'b01000000011001101011100001110111;
		#400 //-5.700688e+25 * -6.3238135e-26 = 3.6050088
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111001010101110101101000001;
		b = 32'b01101010110101010100010011001000;
		correct = 32'b11100010100011100110001110101001;
		#400 //-1.0187564e-05 * 1.28913005e+26 = -1.3133095e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111011100101010011010010100001;
		b = 32'b11011010011001010101010101100111;
		correct = 32'b01010110100001011010100111011011;
		#400 //-0.004553393 * -1.6137918e+16 = 73482285000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111110001000000011100110001;
		b = 32'b11000001011011011010010001000111;
		correct = 32'b11001001101101011111100001110011;
		#400 //100366.38 * -14.852607 = -1490702.4
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111000111011110001001001000100;
		b = 32'b10111010110110111010100110011110;
		correct = 32'b11110100010011010010001100000111;
		#400 //3.8791544e+34 * -0.0016758924 = -6.5010455e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001101100001001001100001010100;
		b = 32'b11101110001110000000010011110100;
		correct = 32'b10111100001111101010000000011010;
		#400 //8.1718e-31 * -1.4237807e+28 = -0.011634851
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010010100110100100000111110101;
		b = 32'b11000000010011001110010011101000;
		correct = 32'b10010011011101101110110011111100;
		#400 //9.735026e-28 * -3.2014713 = -3.1166408e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101110000110111110100010100000;
		b = 32'b00011010111010100010111110011001;
		correct = 32'b01001001100011101001111110011111;
		#400 //1.2062851e+28 * 9.685703e-23 = 1168371.9
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011111010000011101010010000001;
		b = 32'b01010000011000110101100110110111;
		correct = 32'b10110000001011000010001101011100;
		#400 //-4.104512e-20 * 15257230000.0 = -6.2623484e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011011110011011001100000011100;
		b = 32'b01000011000001000000010011001101;
		correct = 32'b10011111010101000000110010010011;
		#400 //-3.4012703e-22 * 132.01875 = -4.4903147e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110000100110001101011101101111;
		b = 32'b11000110111011011100110001001010;
		correct = 32'b01111000000011011111100101101010;
		#400 //-3.784173e+29 * -30438.145 = 1.1518321e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001000011100011100001001000000;
		b = 32'b11010101010111100010110000100100;
		correct = 32'b00011110010100011101000000100011;
		#400 //-7.275164e-34 * -15267573000000.0 = 1.11074095e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110001110001111111011101101011;
		b = 32'b00010001010001010011001010101100;
		correct = 32'b00000011100110100000100011111010;
		#400 //5.8197904e-09 * 1.5556174e-28 = 9.053367e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101101001111001000100111110111;
		b = 32'b01000010101110101100001000001110;
		correct = 32'b10110000100010011000101100101000;
		#400 //-1.0717197e-11 * 93.37901 = -1.0007613e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100100110111011100100011110000;
		b = 32'b10100000000110011001001111000001;
		correct = 32'b00000101100001010000110100011001;
		#400 //-9.6183873e-17 * -1.3008492e-19 = 1.2512071e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110011100001000111011001110011;
		b = 32'b10010000011101010000001101001010;
		correct = 32'b10000100011111011000111000011111;
		#400 //6.168275e-08 * -4.8320264e-29 = -2.9805266e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011111100010011111001011110110;
		b = 32'b00110000010011000110111000111010;
		correct = 32'b01010000010111000101001000000011;
		#400 //1.9880556e+19 * 7.437141e-10 = 14785449000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101101100100100010010101001111;
		b = 32'b10100101110001011100011111011101;
		correct = 32'b01010011111000011101000110011110;
		#400 //-5.6537393e+27 * -3.4309485e-16 = 1939768900000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010111011010100000011111011010;
		b = 32'b10101100000011001111011111010111;
		correct = 32'b10000100000000001101111011011101;
		#400 //7.561939e-25 * -2.0032775e-12 = -1.5148661e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100100111010101010011101110111;
		b = 32'b10001011101001000100011001011001;
		correct = 32'b10110001000101101001001111000100;
		#400 //3.4628842e+22 * -6.327635e-32 = -2.1911868e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001000011110101100011100001011;
		b = 32'b01011010101101011101010101111100;
		correct = 32'b10100011101100100001111111011100;
		#400 //-7.5465612e-34 * 2.559085e+16 = -1.9312292e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100001101011100101000100101110;
		b = 32'b11000001101110110101010010010110;
		correct = 32'b01100011111111110001110111001011;
		#400 //-4.019479e+20 * -23.416302 = 9.412133e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111001100111111101000111000101;
		b = 32'b10000001011111000101010000000011;
		correct = 32'b00111011100111011000011011110001;
		#400 //-1.0372873e+35 * -4.6345366e-38 = 0.004807346
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101000010111000000100110000010;
		b = 32'b11101101011000100111111010110000;
		correct = 32'b11010110010000101010110101001001;
		#400 //1.2214515e-14 * -4.381048e+27 = -53512377000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101101011010010101111110001110;
		b = 32'b01000101010000111011011011001111;
		correct = 32'b01110011001100100110101001110000;
		#400 //4.5140954e+27 * 3131.4255 = 1.4135554e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110101111110110000110010000010;
		b = 32'b11110111110110010110100110101011;
		correct = 32'b01101110010101010011010100111010;
		#400 //-1.8704598e-06 * -8.8193095e+33 = 1.6496164e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101100100001110110010000100100;
		b = 32'b01010000101001010111000101001000;
		correct = 32'b11111101101011101111111011101001;
		#400 //-1.3094231e+27 * 22205317000.0 = -2.9076155e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001011011010010001001100110000;
		b = 32'b01101111011100011000110111111110;
		correct = 32'b10111011010110111110110001010111;
		#400 //-4.4888603e-32 * 7.4757545e+28 = -0.0033557618
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001101001000100101111110010100;
		b = 32'b11000101110110000100101111110001;
		correct = 32'b11010011100010010011000011010000;
		#400 //170260800.0 * -6921.4927 = -1178458900000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000110101001101000000011000010;
		b = 32'b00001111011001001111110011000101;
		correct = 32'b10010110100101001110111100010100;
		#400 //-21312.379 * 1.12899495e-29 = -2.406157e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100110111011100010011110010000;
		b = 32'b00101100001101010010101101001100;
		correct = 32'b10010011101010001000101001000000;
		#400 //-1.6525291e-15 * 2.5745682e-12 = -4.2545487e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001110001000101000101110010010;
		b = 32'b00000100010001100000101111111011;
		correct = 32'b00010010111110110111111100011101;
		#400 //681764000.0 * 2.328029e-36 = 1.5871663e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101000010111101100100001111101;
		b = 32'b01000101000000111111010111101011;
		correct = 32'b11101101111001011010110100110101;
		#400 //-4.208255e+24 * 2111.3699 = -8.885183e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110000001000101111001011110010;
		b = 32'b00110000010001011010010000000000;
		correct = 32'b01100000111110111001101010110000;
		#400 //2.017211e+29 * 7.190124e-10 = 1.4503997e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000001100000001101001001001010;
		b = 32'b11001001011100001000100010010111;
		correct = 32'b00001011011100100001001111000010;
		#400 //-4.7321524e-38 * -985225.44 = 4.662237e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000010000001001111111000101011;
		b = 32'b01001101110001010100011100100011;
		correct = 32'b01010000010011001111100100011000;
		#400 //33.24821 * 413721700.0 = 13755507000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011000111110111011101111000101;
		b = 32'b01111100010001011000101000110010;
		correct = 32'b11010101110000100011111101100011;
		#400 //-6.507158e-24 * 4.1027417e+36 = -26697187000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110001010111111111010101100010;
		b = 32'b00011101011110111110100100010100;
		correct = 32'b00001111010111000110000101111111;
		#400 //3.2590255e-09 * 3.3340072e-21 = 1.08656145e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101010100011110110111111000010;
		b = 32'b10110010111001110111111001100010;
		correct = 32'b00011110000000011011010010101000;
		#400 //-2.547945e-13 * -2.6949412e-08 = 6.866562e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011010000111001111111000001000;
		b = 32'b01100100001110101101011100100010;
		correct = 32'b00111110111001010010100100000000;
		#400 //3.246525e-23 * 1.3786385e+22 = 0.44757843
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011000100011000111111110111100;
		b = 32'b10111110101000011000111101110100;
		correct = 32'b11010111101100010101011000100000;
		#400 //1235842000000000.0 * -0.3155476 = -389966920000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110110011101001011100100100100;
		b = 32'b00010100001001100100100101111100;
		correct = 32'b11001011000111101111011001001101;
		#400 //-1.2408941e+33 * 8.3953505e-27 = -10417741.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100011101100011110010111011101;
		b = 32'b01101001010111000010010110101101;
		correct = 32'b01001101100110001111101110111000;
		#400 //1.928773e-17 * 1.663385e+25 = 320829200.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101000000011110001111100000010;
		b = 32'b10101000100100011000001101100100;
		correct = 32'b01010001001000101011010000001010;
		#400 //-2.7034816e+24 * -1.6155215e-14 = 43675330000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010001110011110001101011000111;
		b = 32'b00011110010111101010110111100001;
		correct = 32'b00110000101101000010010111100100;
		#400 //111188435000.0 * 1.17885395e-20 = 1.3107493e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001011110111011001100000000011;
		b = 32'b11111000111010001100100000000101;
		correct = 32'b11000101010010010111111011100110;
		#400 //8.5354825e-32 * -3.777093e+34 = -3223.9312
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101110000010110010110010111101;
		b = 32'b00111101001000001011100000101011;
		correct = 32'b01101011101011101100000000101011;
		#400 //1.0768125e+28 * 0.039238136 = 4.2252116e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011101010101110100110100111101;
		b = 32'b11011000101010001000010100100110;
		correct = 32'b01110110100011011011101010101011;
		#400 //-9.696327e+17 * -1482318600000000.0 = 1.4373046e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011100101110100100110101001111;
		b = 32'b10010010010000011101011100000111;
		correct = 32'b10101111100011010001000011000101;
		#400 //4.1951478e+17 * -6.1165104e-28 = -2.5659666e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001110010000001011001011101011;
		b = 32'b00101100011011001100100111000001;
		correct = 32'b00111011001100100011110011001110;
		#400 //808237760.0 * 3.3649613e-12 = 0.0027196887
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011000101001111101110000001110;
		b = 32'b00111010100110000111000010101100;
		correct = 32'b00010011110001111110100100010011;
		#400 //4.3390687e-24 * 0.0011630259 = 5.046449e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010001001100000010001011011111;
		b = 32'b00110101110000101011011101011011;
		correct = 32'b11000111100001011111100010010101;
		#400 //-47281205000.0 * 1.450749e-06 = -68593.164
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101000111101100100101001100101;
		b = 32'b10101101000100100001100011001100;
		correct = 32'b11010110100011001000111001001001;
		#400 //9.304596e+24 * -8.304645e-12 = -77271370000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101011100000010000101100101011;
		b = 32'b10111110000100000000010000001001;
		correct = 32'b11101010000100010011000010100010;
		#400 //3.1200834e+26 * -0.1406404 = -4.3880976e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001001001000101101001011100000;
		b = 32'b11011001100100001000110010110111;
		correct = 32'b11100011001101111110000000111011;
		#400 //666926.0 * -5085889300000000.0 = -3.3919117e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110010011010100111100111001000;
		b = 32'b10111010000000100110001011000111;
		correct = 32'b10101100111011101101100010100001;
		#400 //1.36482825e-08 * -0.00049738254 = -6.7884175e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100110011101110100001100101000;
		b = 32'b11001011100100110011001001110110;
		correct = 32'b11110010100011100010110001001101;
		#400 //2.9191583e+23 * -19293420.0 = -5.632055e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010110100011001110111100101000;
		b = 32'b01110111010000101111100010001101;
		correct = 32'b01001110010101101010110000100011;
		#400 //2.2769149e-25 * 3.9544797e+33 = 900401340.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101101100010100100011101011111;
		b = 32'b11000001000010001010101011100101;
		correct = 32'b11101111000100111010010001110011;
		#400 //5.349402e+27 * -8.541722 = -4.5693103e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111101010100011110101101010101;
		b = 32'b11010000111101001101000011111010;
		correct = 32'b11001110110010001011111110101001;
		#400 //0.05124982 * -32858690000.0 = -1684001900.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011101111111010100001011111000;
		b = 32'b11011010110111100110010000001100;
		correct = 32'b11111001010111000000001100001101;
		#400 //2.2811777e+18 * -3.1298724e+16 = -7.139795e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010010010000100111110101000000;
		b = 32'b10011000111111101101000011110010;
		correct = 32'b00101011110000011001011100000011;
		#400 //-208831250000.0 * -6.586844e-24 = 1.3755389e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101011111101110100000011011110;
		b = 32'b10100000010010010110010011111101;
		correct = 32'b10001100110000101000001101111000;
		#400 //1.756841e-12 * -1.7058776e-19 = -2.9969558e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000001001010010101001001100000;
		b = 32'b00011100100011101000101101001100;
		correct = 32'b10011110001111001000111110100110;
		#400 //-10.582611 * 9.432779e-22 = -9.982343e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001100010001110000111100001100;
		b = 32'b11000101110010011010011010011001;
		correct = 32'b11010010100111001100110001011011;
		#400 //52182064.0 * -6452.8247 = -336721700000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110011000101110100011000101011;
		b = 32'b11100111111100100111110100111001;
		correct = 32'b01011011100011110100101001010100;
		#400 //-3.5221245e-08 * -2.2902453e+24 = 8.066529e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101010111000100110100000001111;
		b = 32'b01000110000111011011010001001000;
		correct = 32'b00110001100010110111100101000010;
		#400 //4.021787e-13 * 10093.07 = 4.059218e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111011111101010011010000010110;
		b = 32'b10111001000100110100110000100010;
		correct = 32'b01110101100011010001010111010101;
		#400 //-2.5463383e+36 * -0.00014047374 = 3.576937e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010011010101101010101110011100;
		b = 32'b01011010001101111001011100110100;
		correct = 32'b10101110000110011111001101110111;
		#400 //-2.7095207e-27 * 1.2919043e+16 = -3.5004413e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010011100110011000100001101000;
		b = 32'b11001100111011000101000010011101;
		correct = 32'b00100001000011011011101000011001;
		#400 //-3.8757137e-27 * -123897064.0 = 4.8018956e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111001110011011000111001101010;
		b = 32'b01000100110000010100110010011110;
		correct = 32'b10111111000110110011010111100011;
		#400 //-0.00039206754 * 1546.3943 = -0.606291
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000000101011101010111010101010;
		b = 32'b01010000001100001110000000111000;
		correct = 32'b00010001011100010110001000101000;
		#400 //1.6042034e-38 * 11869938000.0 = 1.9041795e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011110000011110010100001111111;
		b = 32'b00101101110001111100010111001001;
		correct = 32'b10001100010111110110111000101011;
		#400 //-7.578731e-21 * 2.2711515e-11 = -1.7212448e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111000001101000011010001001000;
		b = 32'b00011101000100001001100110010011;
		correct = 32'b00010101110010111001001100000110;
		#400 //4.2964035e-05 * 1.9137637e-21 = 8.222301e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001111011011001001001001101000;
		b = 32'b00011101000001011101111110001010;
		correct = 32'b10101100111101110110110101000110;
		#400 //-3969017900.0 * 1.771797e-21 = -7.032294e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100001010111010010110100000101;
		b = 32'b00100110000010001001001010001100;
		correct = 32'b01000111111010111111110100001111;
		#400 //2.549984e+20 * 4.7383087e-16 = 120826.12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100101111010001100101100010101;
		b = 32'b01100011000111110111001010111101;
		correct = 32'b01001001100100001111111001111000;
		#400 //4.0383198e-16 * 2.9413e+21 = 1187791.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110110010110110100111011111100;
		b = 32'b10010101100101100001000001110111;
		correct = 32'b10001100100000001000111001100011;
		#400 //3.2679518e-06 * -6.0610494e-26 = -1.9807219e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110010000011100110111110010010;
		b = 32'b01001110000000111100010011011000;
		correct = 32'b11000000100100101010000100111011;
		#400 //-8.290856e-09 * 552678900.0 = -4.5821815
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001100100111000100100100100101;
		b = 32'b01101111101100101010100000000101;
		correct = 32'b11111100110110100010001011011110;
		#400 //-81938730.0 * 1.1058291e+29 = -9.061023e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010110111110100101101110111010;
		b = 32'b01011010001111011010001000101111;
		correct = 32'b10110001101110010111010001010100;
		#400 //-4.0447566e-25 * 1.3344273e+16 = -5.3974336e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100011001000110011011100000001;
		b = 32'b11011000100100010100101010111001;
		correct = 32'b10111100001110010100001110010111;
		#400 //8.847895e-18 * -1278001000000000.0 = -0.011307619
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001011001111001010011001010001;
		b = 32'b11101100000101011101001101100111;
		correct = 32'b10110111110111001101000100101100;
		#400 //3.6332606e-32 * -7.245131e+26 = -2.6323447e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011100101011111000010000111000;
		b = 32'b10101000100000000001110110000111;
		correct = 32'b00000101101011111010110010110101;
		#400 //-1.1614706e-21 * -1.422366e-14 = 1.6520363e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100010100001010000000111000001;
		b = 32'b01001010010101111110101011010001;
		correct = 32'b00101101011000000101110011110011;
		#400 //3.605158e-18 * 3537588.2 = 1.2753565e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001111110110111011110100011000;
		b = 32'b01000101000110010011100010111011;
		correct = 32'b11010101100000111000010010110101;
		#400 //-7373205500.0 * 2451.5457 = -18075750000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100100101111010100101100010101;
		b = 32'b00100101111000011101111110101110;
		correct = 32'b01001011001001110000010001100011;
		#400 //2.793476e+22 * 3.918285e-16 = 10945635.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100010101110100010100010111011;
		b = 32'b11110111110110000010101001010011;
		correct = 32'b01011011000111010011000100100101;
		#400 //-5.0458526e-18 * -8.7687075e+33 = 4.4245606e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100001000010101011110101111110;
		b = 32'b11010110011010101001010101111100;
		correct = 32'b10110111111111100100010001110001;
		#400 //4.700701e-19 * -64481938000000.0 = -3.031103e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110100111011010110101011001;
		b = 32'b11101000001100011100110001100001;
		correct = 32'b11100111010110110000010101111001;
		#400 //0.30796316 * -3.358516e+24 = -1.0342992e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000011100011110100010110100100;
		b = 32'b11010001110001101000111111011001;
		correct = 32'b10010101110111100100000010111100;
		#400 //8.420773e-37 * -106602110000.0 = -8.976722e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001111101100000001010010111001;
		b = 32'b00110111111000000110100010011010;
		correct = 32'b11001000000110100101101000010100;
		#400 //-5908296000.0 * 2.675159e-05 = -158056.31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110000000010111111001001100000;
		b = 32'b00010001100110110110100001101010;
		correct = 32'b00000010001010011110100110101001;
		#400 //5.091234e-10 * 2.4519038e-28 = 1.2483216e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011010110111101101000000111011;
		b = 32'b11011001011100001111111110110111;
		correct = 32'b00110100110100011100000111001000;
		#400 //-9.215346e-23 * -4239697200000000.0 = 3.9070278e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001011100111111010011000010110;
		b = 32'b10000110111111011110111001110100;
		correct = 32'b10010011000111100101101111011000;
		#400 //20925484.0 * -9.55184e-35 = -1.9987686e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001010110000110100000110011010;
		b = 32'b10000110100001110101000010010100;
		correct = 32'b00010001110011100110101000011011;
		#400 //-6398157.0 * -5.0899755e-35 = 3.2566462e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011110111101001010111101101010;
		b = 32'b01011011001110100100011101100111;
		correct = 32'b11111010101100100000101110110010;
		#400 //-8.815714e+18 * 5.2432853e+16 = -4.6223302e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011011110011100111111011000010;
		b = 32'b01100100010001010000000011100101;
		correct = 32'b01000000100111101110100001000100;
		#400 //3.4161757e-22 * 1.4536292e+22 = 4.9658527
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111000010110100011001000000100;
		b = 32'b00011110111111101001011101000111;
		correct = 32'b10010111110110001111111010010000;
		#400 //-5.202183e-05 * 2.6955863e-20 = -1.4022933e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100111100110000111011111101101;
		b = 32'b11000000101000001111111011111100;
		correct = 32'b01101000101111111100010110100010;
		#400 //-1.4400239e+24 * -5.031126 = 7.2449414e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001110101010010001001000001110;
		b = 32'b01001011101110011000100111101100;
		correct = 32'b10011010111101010001001001000101;
		#400 //-4.1679103e-30 * 24318936.0 = -1.0135914e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101010110101100001000011010100;
		b = 32'b00100011011100111011010001111010;
		correct = 32'b00001110110010111100100011100011;
		#400 //3.8025713e-13 * 1.3211274e-17 = 5.023681e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101111001011100010111011111001;
		b = 32'b01000100001100101101011110000101;
		correct = 32'b10110011111100110101111010011010;
		#400 //-1.5841896e-10 * 715.3675 = -1.1332777e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110111011011000110010111011011;
		b = 32'b11111101101000010001110100111011;
		correct = 32'b11110101100101001100011100001101;
		#400 //1.4090411e-05 * -2.6769685e+37 = -3.771959e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111001101110010001110110011010;
		b = 32'b10010000011110110110110000010101;
		correct = 32'b11001010101101011100111000101110;
		#400 //1.2014691e+35 * -4.9584285e-29 = -5957399.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000111110100110110001110011101;
		b = 32'b11000010001101111100100111110001;
		correct = 32'b01001010100101111100001011110101;
		#400 //-108231.23 * -45.94721 = 4972922.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000001100111001010100110101100;
		b = 32'b01100101001101000000111011000101;
		correct = 32'b00100111010111000110000010101110;
		#400 //5.7548817e-38 * 5.314365e+22 = 3.0583543e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101001111100011110110100001001;
		b = 32'b10001011000000001101111101010111;
		correct = 32'b00110101011100111001001100101000;
		#400 //-3.6558811e+25 * -2.4819926e-32 = 9.0738695e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100110011101001010111100010100;
		b = 32'b11011111010011100111110110001111;
		correct = 32'b11000110010001010101110011100100;
		#400 //8.489178e-16 * -1.4879206e+19 = -12631.223
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111000000110110001000010100010;
		b = 32'b11000101011100110101001101110101;
		correct = 32'b01111110000100110110001101010111;
		#400 //-1.2580365e+34 * -3893.216 = 4.897808e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011000001001101000011111101100;
		b = 32'b01101101000101000011010001111001;
		correct = 32'b11000101110000001101000101101110;
		#400 //-2.152362e-24 * 2.866701e+27 = -6170.1787
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111100011011010010111110110111;
		b = 32'b00010011110100001000110001011001;
		correct = 32'b01010000110000010011100011001101;
		#400 //4.9261685e+36 * 5.2644975e-27 = 25933801000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010110001001101001000100110000;
		b = 32'b00101101111110001101101111100011;
		correct = 32'b11000100101000011110101110111000;
		#400 //-45785626000000.0 * 2.8291985e-11 = -1295.3662
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101100110111100101011000000100;
		b = 32'b00011010000111000001001011000011;
		correct = 32'b01000111100001111000110010110110;
		#400 //2.1503018e+27 * 3.22752e-23 = 69401.42
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101001000101101100001110010001;
		b = 32'b11010001110010111110000011111101;
		correct = 32'b00111011011100000010001100101000;
		#400 //-3.3476318e-14 * -109456630000.0 = 0.0036642049
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111110101111000001111011111111;
		b = 32'b00110001110111101000010001101001;
		correct = 32'b11110001001000111000010000101110;
		#400 //-1.250279e+38 * 6.4761037e-09 = -8.096936e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101111110011100011010000111101;
		b = 32'b00101110101011000111000100110101;
		correct = 32'b01011111000010101110011001001001;
		#400 //1.2763413e+29 * 7.841764e-11 = 1.0008767e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100101010000001001010100011111;
		b = 32'b00101000000010111111010001010110;
		correct = 32'b00001101110100101001000110001101;
		#400 //1.670387e-16 * 7.769032e-15 = 1.2977289e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011100100110111011010001100111;
		b = 32'b01011011100001110101000011000101;
		correct = 32'b10111000101001001001101010000101;
		#400 //-1.0303673e-21 * 7.617586e+16 = -7.848911e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010001011000110011101001110011;
		b = 32'b01110000110010111001011110110000;
		correct = 32'b11000010101101001011010111111101;
		#400 //-1.7925154e-28 * 5.040707e+29 = -90.355446
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010001111001000011101010000011;
		b = 32'b11001101010100110100111111001110;
		correct = 32'b11011111101111000110001101100000;
		#400 //122529276000.0 * -221576420.0 = -2.7149599e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101011110110101000001000011011;
		b = 32'b10010111100011111111011111001010;
		correct = 32'b11000011111101011100010001011010;
		#400 //5.2832047e+26 * -9.303709e-25 = -491.534
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011011001010100101110110001000;
		b = 32'b01010010011101001000101111110101;
		correct = 32'b00101110001000101011111001001001;
		#400 //1.4092292e-22 * 262580030000.0 = 3.7003543e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100000101100011011010000101100;
		b = 32'b10101011110110011010110011001011;
		correct = 32'b00001101000101110001100110101011;
		#400 //-3.0104194e-19 * -1.5466737e-12 = 4.6561364e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000110100001011001001101010001;
		b = 32'b00011010110000011110110100100100;
		correct = 32'b10100001110010100101111110011000;
		#400 //-17097.658 * 8.020605e-23 = -1.3713356e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111011011000010100110010011110;
		b = 32'b10111010001111010000100011111011;
		correct = 32'b01110110001001100101110101111000;
		#400 //-1.1698208e+36 * -0.0007211116 = 8.435713e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101111001110101011011100011100;
		b = 32'b00101001011100101001010101000100;
		correct = 32'b10011001001100001110110111110111;
		#400 //-1.6981655e-10 * 5.386426e-14 = -9.147043e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001111010111100001101011010000;
		b = 32'b01011000010100100111100001011000;
		correct = 32'b11101000001101101001101001101000;
		#400 //-3726299100.0 * 925657260000000.0 = -3.449276e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111000100111011110010101010;
		b = 32'b01010110110011010111011101001110;
		correct = 32'b11001110011011010010010111011100;
		#400 //-8.80581e-06 * 112956150000000.0 = -994670340.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001001110111010100010010010001;
		b = 32'b11101110111010000100000011110101;
		correct = 32'b11111001010010001011111001001000;
		#400 //1812626.1 * -3.5939525e+28 = -6.514492e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001100011000011000010110010011;
		b = 32'b11010010010100000000011100011011;
		correct = 32'b10011111001101110100001011001010;
		#400 //1.7373566e-31 * -223368100000.0 = -3.8807004e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101001010010111010101100010111;
		b = 32'b11000110011011110110111001011010;
		correct = 32'b10110000001111100111110010000110;
		#400 //4.522345e-14 * -15323.588 = -6.9298556e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110100111000010100110111111100;
		b = 32'b10111011100110100001110101100001;
		correct = 32'b00110001000001111010001011000101;
		#400 //-4.1966257e-07 * -0.0047032093 = 1.973761e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000101010011000011101000000000;
		b = 32'b11110110100011110110010011110111;
		correct = 32'b11111100011001001100100111100011;
		#400 //3267.625 * -1.4541919e+33 = -4.7517537e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111100100010110111000110011010;
		b = 32'b11111110101000000000110011111101;
		correct = 32'b11111011101011100101110000100111;
		#400 //0.017021943 * -1.0637196e+38 = -1.8106574e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101111011010111000000000001101;
		b = 32'b11101110100110110110100010111100;
		correct = 32'b11011110100011101111011011100001;
		#400 //2.1418618e-10 * -2.4048396e+28 = -5.1508343e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110011100001101101010100011100;
		b = 32'b01010110111100011000010111101111;
		correct = 32'b01001010111111100110101001010100;
		#400 //6.2786256e-08 * 132778770000000.0 = 8336682.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011100001010011000101011000000;
		b = 32'b01100000100000111101011100010000;
		correct = 32'b11111101001011101010000011011101;
		#400 //-1.9088731e+17 * 7.600064e+19 = -1.4507558e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011101110100100000100000011110;
		b = 32'b00111011010000000011110000011001;
		correct = 32'b10011001100111011011011101100101;
		#400 //-5.559493e-21 * 0.0029332696 = -1.6307492e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000101110110101111011011101111;
		b = 32'b11010011011011011111001011001111;
		correct = 32'b01011001110010111000011001001010;
		#400 //-7006.8667 * -1021980900000.0 = 7160884000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000010011111111001110011111111;
		b = 32'b10000000000001110100100100011000;
		correct = 32'b10000001011010001100100011010111;
		#400 //63.903316 * -6.6907e-40 = -4.2755766e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111011010111110000011101100010;
		b = 32'b10011011010110010010110100001011;
		correct = 32'b10010111001111010011010010000000;
		#400 //0.00340315 * -1.7964373e-22 = -6.113546e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011110010111101000110001010;
		b = 32'b10010010111001010011010011000110;
		correct = 32'b00011111001101100111110001110101;
		#400 //-26714900.0 * -1.4464941e-27 = 3.8642948e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110000100011111000111101011111;
		b = 32'b11011111010011001011001001100100;
		correct = 32'b11010000011001011001010010010011;
		#400 //1.0445368e-09 * -1.4749962e+19 = -15406878000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101110110101111111101010110110;
		b = 32'b10001000011101110011010010000101;
		correct = 32'b00110111110100001000111100110101;
		#400 //-3.3421184e+28 * -7.4390595e-34 = 2.4862218e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100000110101111101100001000110;
		b = 32'b11100111111011100110111111100100;
		correct = 32'b01001001010010010000100101101000;
		#400 //-3.6565534e-19 * -2.2519745e+24 = 823446.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110010011011010000101101100111;
		b = 32'b10110110011111000011010010001000;
		correct = 32'b11101001011010011000011111011110;
		#400 //4.6951508e+30 * -3.7581503e-06 = -1.7645083e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100011101101111111100101111110;
		b = 32'b00010011100101111101101101001111;
		correct = 32'b00110111110110100100001110001001;
		#400 //6.787464e+21 * 3.8334014e-27 = 2.6019074e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011011110101101100110110110010;
		b = 32'b00001101011100100101110101110101;
		correct = 32'b00101001110010110101110011011101;
		#400 //1.2092362e+17 * 7.46845e-31 = 9.03112e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000111111010101100011011111100;
		b = 32'b01101011111010010001101010111110;
		correct = 32'b10110100010101011100011110100010;
		#400 //-3.532536e-34 * 5.63612e+26 = -1.9909797e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111001100101101000110000000;
		b = 32'b00111010000110000100101000001011;
		correct = 32'b01000001110101001100000000111000;
		#400 //45777.5 * 0.0005809373 = 26.593857
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001011001110111011101011101100;
		b = 32'b00111100011001011101001111011010;
		correct = 32'b10001000001010001000100110010000;
		#400 //-3.6155514e-32 * 0.01402756 = -5.0717365e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000001101100110011111100000001;
		b = 32'b00100001111010000011011001001111;
		correct = 32'b00100100001000101001011100100000;
		#400 //22.405764 * 1.5735307e-18 = 3.5256158e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001110011010000101001000100100;
		b = 32'b10110110011101011100100101111011;
		correct = 32'b01000101010111110000110101110101;
		#400 //-974424300.0 * -3.6625122e-06 = 3568.841
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010110101111010110000110101001;
		b = 32'b11010100101100010000100100101010;
		correct = 32'b10101100000000101111011101001101;
		#400 //3.059623e-25 * -6082903700000.0 = -1.861139e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010100100111001011001011111101;
		b = 32'b10110101000111101010000100100111;
		correct = 32'b10001010010000100011001000111001;
		#400 //1.5822573e-26 * -5.9094094e-07 = -9.350206e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000101101011011101101011001010;
		b = 32'b00101110100110000111001110001000;
		correct = 32'b00110100110011110001000010111011;
		#400 //5563.3486 * 6.932682e-11 = 3.8568928e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101111000000000001001010101011;
		b = 32'b11011001111001000110001000010001;
		correct = 32'b11001001011001001000001101100000;
		#400 //1.1648164e-10 * -8035515000000000.0 = -935990.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010111000010100000110000001110;
		b = 32'b11001010101011101110101100011011;
		correct = 32'b11100010001111001010010111110010;
		#400 //151784380000000.0 * -5731725.5 = -8.699864e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111011101001111111111001001010;
		b = 32'b00000110000010100100011010110100;
		correct = 32'b01000010001101010111101011110011;
		#400 //1.7445423e+36 * 2.600686e-35 = 45.370068
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010011001101111010110001100100;
		b = 32'b00101011010101111010111100101010;
		correct = 32'b00111111000110101011111101110101;
		#400 //788871250000.0 * 7.6626433e-13 = 0.6044839
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001001000000110101100110000001;
		b = 32'b01010100011001110111110100101001;
		correct = 32'b10011101111011011000101111110110;
		#400 //-1.5810636e-33 * 3976949100000.0 = -6.2878094e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010100011001101111110100001011;
		b = 32'b10100001010110001010010010010110;
		correct = 32'b10110110010000110111101000000011;
		#400 //3968351300000.0 * -7.3401474e-19 = -2.9128284e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111011110000000110010011101;
		b = 32'b11011100101111111111011011000100;
		correct = 32'b01010100101110100000000010000011;
		#400 //-1.4784889e-05 * -4.3226434e+17 = 6390980000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011011011010111011111001011110;
		b = 32'b10110111111000100010011101111000;
		correct = 32'b01010011110100000100001001100111;
		#400 //-6.635593e+16 * -2.6959679e-05 = 1788934500000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100010011110010101101100000111;
		b = 32'b00110001100010110010111100100110;
		correct = 32'b01010100100001111001001001011010;
		#400 //1.1499496e+21 * 4.0507926e-09 = 4658207700000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110000100101100100111011110000;
		b = 32'b01010001011101110011111011001001;
		correct = 32'b01000010100100010010101100000111;
		#400 //1.0936372e-09 * 66369393000.0 = 72.58404
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011110001001100111111010000001;
		b = 32'b00010111010011101100101110010101;
		correct = 32'b00110110000001100111111000110011;
		#400 //2.999292e+18 * 6.6819147e-25 = 2.0041014e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101000011101111111110110001010;
		b = 32'b00100001011001100101011111101001;
		correct = 32'b11001010010111110010001011110011;
		#400 //-4.684406e+24 * 7.804338e-19 = -3655868.8
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011010000011110110001110111010;
		b = 32'b10010101000111001010011100010110;
		correct = 32'b10101111101011110111110010110111;
		#400 //1.0090143e+16 * -3.1635757e-26 = -3.192093e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111000111000111011000011011000;
		b = 32'b10111110110111001101100100100111;
		correct = 32'b00111000010001000110110100011101;
		#400 //-0.00010857143 * -0.43134424 = 4.683166e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111100010110111110101100100100;
		b = 32'b10111100111001100110000110010101;
		correct = 32'b11111001110001011110100100010110;
		#400 //4.567529e+36 * -0.028122703 = -1.2845125e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110111111101010100101101111110;
		b = 32'b10100000000010000011110101001010;
		correct = 32'b11011000100000101000101011010101;
		#400 //9.950343e+33 * -1.1539927e-19 = -1148262300000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101100000001100011100010110010;
		b = 32'b01100011001001110010100110111011;
		correct = 32'b01001111101011110100100110111010;
		#400 //1.9074018e-12 * 3.0836133e+21 = 5881689000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011100010010000110111101111111;
		b = 32'b00101100110000000111000110100111;
		correct = 32'b00001001100101101010110010011011;
		#400 //6.6318554e-22 * 5.469586e-12 = 3.6273504e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111000110011010010100001111000;
		b = 32'b00000011001011110001100001101000;
		correct = 32'b10111100100011000101001000111001;
		#400 //-3.3288802e+34 * 5.1455895e-37 = -0.01712905
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001101001011010000111111111100;
		b = 32'b01011101101110011001011100111001;
		correct = 32'b01101011011110101110110110010000;
		#400 //181469120.0 * 1.6716525e+18 = 3.0335331e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001111001001011100111100101111;
		b = 32'b01011010110100000111010001101001;
		correct = 32'b00101010100001110000001110111100;
		#400 //8.17503e-30 * 2.9337395e+16 = 2.3983409e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000101101001110101011111111;
		b = 32'b10100011110001111111101110111101;
		correct = 32'b00010101000011010101010010010100;
		#400 //-1.3163514e-09 * -2.1682239e-17 = 2.8541444e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100100011111101100100101101010;
		b = 32'b11011011110001010000011001100111;
		correct = 32'b01000000110001000001011101011110;
		#400 //-5.5248075e-17 * -1.1091522e+17 = 6.1278524
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110101010101001001101000001011;
		b = 32'b10011111000010000100110000110010;
		correct = 32'b01010100111000100110001000111010;
		#400 //-2.6950471e+32 * -2.8862147e-20 = 7778484600000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111000001000010000110010010001;
		b = 32'b10111111111100000110011110111111;
		correct = 32'b00111000100101110011110100001100;
		#400 //-3.8397095e-05 * -1.8781661 = 7.211612e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100011110001110101100010101101;
		b = 32'b11000101110000000110111100110100;
		correct = 32'b10101010000101011101100100011010;
		#400 //2.1613179e-17 * -6157.9004 = -1.3309181e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011101010010000011001011111100;
		b = 32'b10001011000001101010100111001001;
		correct = 32'b00101000110100101001111011101110;
		#400 //-9.0161685e+17 * -2.5935193e-32 = 2.3383608e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000010111000110010101110110001;
		b = 32'b10001111101110111101111101000000;
		correct = 32'b00010011001001101011011100000110;
		#400 //-113.585335 * -1.8525616e-29 = 2.1042383e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100000101101010101101111101110;
		b = 32'b11010111010101010011101011010011;
		correct = 32'b11111000100101110000111100101001;
		#400 //1.045464e+20 * -234448620000000.0 = -2.451076e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110100010100000110010001001010;
		b = 32'b11111111000110011011111111000111;
		correct = 32'b01110011111110100101000000011010;
		#400 //-1.9407995e-07 * -2.0436765e+38 = 3.9663662e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101111001111001110101011011010;
		b = 32'b10101111110100110011000010111001;
		correct = 32'b10011111100110111101100110000110;
		#400 //1.7181936e-10 * -3.8415296e-10 = -6.6004916e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011111000101000011000111100100;
		b = 32'b00000111010000100101010001001010;
		correct = 32'b10100110111000001111110100110100;
		#400 //-1.0678567e+19 * 1.4619708e-34 = -1.5611753e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110110010101111100000001101000;
		b = 32'b00111100011001100010101101100100;
		correct = 32'b01110011010000011111101101101111;
		#400 //1.0939905e+33 * 0.014048431 = 1.536885e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110110110011100111111000011110;
		b = 32'b10101000000110100011111100101101;
		correct = 32'b10011111011110001101010110100111;
		#400 //6.1539604e-06 * -8.562416e-15 = -5.2692772e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100011011000111001010110011100;
		b = 32'b01111000110101100001000001010100;
		correct = 32'b01011100101111100100110110010100;
		#400 //1.2337376e-17 * 3.4733834e+34 = 4.2852435e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110100111110011011001010101001;
		b = 32'b10110111101101000100000000111111;
		correct = 32'b11101101001011111101000001001001;
		#400 //1.5826484e+32 * -2.1487589e-05 = -3.40073e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001011101111010000101001011010;
		b = 32'b11001110100000110011010010010100;
		correct = 32'b10011010110000011100011000111111;
		#400 //7.281573e-32 * -1100630500.0 = -8.014321e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000010111010111010110001101100;
		b = 32'b00110001101100100000100000001011;
		correct = 32'b00110101001000111110010101001011;
		#400 //117.83676 * 5.181396e-09 = 6.1055897e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111101101001111111001100000010;
		b = 32'b00110110111101110110010011011110;
		correct = 32'b11110101001000100100110110100011;
		#400 //-2.7905355e+37 * 7.372916e-06 = -2.0574384e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010011101110100101001001000000;
		b = 32'b01011010101100010001100000100101;
		correct = 32'b00101111000000001110010001110001;
		#400 //4.7034106e-27 * 2.492381e+16 = 1.1722691e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000011111110101011100110001010;
		b = 32'b01110010000100110100001011111010;
		correct = 32'b01110110100100000011101000100011;
		#400 //501.44952 * 2.916817e+30 = 1.4626365e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110100100101101000111100010010;
		b = 32'b10001110011100011101000001001001;
		correct = 32'b10000011100011100011011100101111;
		#400 //2.8043775e-07 * -2.980583e-30 = -8.358679e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011101010111000001101001011001;
		b = 32'b10010011100011110100010100111010;
		correct = 32'b00110001011101100101110001111001;
		#400 //-9.912554e+17 * -3.6166538e-27 = 3.5850276e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111110111110100100111000110001;
		b = 32'b11001001001110100100111111101011;
		correct = 32'b01001000101101100010101011110100;
		#400 //-0.4888778 * -763134.7 = 373079.62
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100111011010100100111110110110;
		b = 32'b10011010000101011001110000111011;
		correct = 32'b00000010000010001110111101100100;
		#400 //-3.2517235e-15 * -3.093868e-23 = 1.0060404e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100110000010011111101100101011;
		b = 32'b11000001011011001011001010001011;
		correct = 32'b11100111111111110010011110001110;
		#400 //1.6289936e+23 * -14.79359 = -2.4098662e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101100110001011100000110111000;
		b = 32'b11010111100101000111110000100001;
		correct = 32'b01000100111001010110011111000011;
		#400 //-5.620584e-12 * -326521700000000.0 = 1835.2426
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001001110001101001111010000011;
		b = 32'b00100101110010001011111101011011;
		correct = 32'b00110000000110111100000001001101;
		#400 //1627088.4 * 3.4824137e-16 = 5.666195e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011000000101001111000000101111;
		b = 32'b01111110110111001111100011100100;
		correct = 32'b11010111100000001000111100110110;
		#400 //-1.9249813e-24 * 1.4686124e+38 = -282705150000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100010111001011010011100101001;
		b = 32'b01011010010101101100110000100001;
		correct = 32'b00111101110000001011000011011011;
		#400 //6.2247562e-18 * 1.5115022e+16 = 0.094087325
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111111010101000001000111111001;
		b = 32'b11110111101110111001101101100010;
		correct = 32'b11110111100110110110100111011001;
		#400 //0.82839924 * -7.6102426e+33 = -6.304319e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111011001000100101010010001100;
		b = 32'b00110001000000010000011000001101;
		correct = 32'b00101100101000111010000011100010;
		#400 //0.0024769632 * 1.877541e-09 = 4.6506002e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100011001000101101001001000010;
		b = 32'b11000000100001110101100111001110;
		correct = 32'b10100100001011000010101111111110;
		#400 //8.8265614e-18 * -4.2297125 = -3.7333818e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001001000110111101011110100110;
		b = 32'b11100001000110010001110001110100;
		correct = 32'b11101010101110100110101001101001;
		#400 //638330.4 * -1.7652513e+20 = -1.12681355e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110101001110100101100001100101;
		b = 32'b00010010111100000111110110100001;
		correct = 32'b01001000101011110000111001010001;
		#400 //2.3622072e+32 * 1.5177099e-27 = 358514.53
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100101110011101001000010000011;
		b = 32'b01010101010101001000000010011011;
		correct = 32'b00111011101010110111011101110010;
		#400 //3.5833229e-16 * 14603051000000.0 = 0.005232745
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011100010100001001011001111101;
		b = 32'b00110011000000111000100001101000;
		correct = 32'b01001111110101100101100001001101;
		#400 //2.3484904e+17 * 3.0624875e-08 = 7192222000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110001111011000000100101111011;
		b = 32'b00110001100010000111010011100111;
		correct = 32'b10100011111110111010000110100101;
		#400 //-6.869582e-09 * 3.971411e-09 = -2.7281934e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101011110101011111000001100000;
		b = 32'b00011110001001110000011010101001;
		correct = 32'b00001010100010111001010101011111;
		#400 //1.5201278e-12 * 8.842284e-21 = 1.34414e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010000100110000110001100110101;
		b = 32'b10000100011101110000111000000011;
		correct = 32'b00010101100100110001000000001111;
		#400 //-20453108000.0 * -2.9041144e-36 = 5.9398163e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110011110001010111101101000;
		b = 32'b01110000001101100010101000111000;
		correct = 32'b11100111001100001111010110110111;
		#400 //-3.705698e-06 * 2.2550924e+29 = -8.3566914e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110010111001110001101111000;
		b = 32'b00100110000110100100100110000001;
		correct = 32'b00100101000001010010000001000010;
		#400 //0.21571147 * 5.35291e-16 = 1.154684e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010001001010010010000111101;
		b = 32'b11111100000101101001011110001111;
		correct = 32'b01110110110000100100101000000001;
		#400 //-0.00062996504 * -3.127674e+36 = 1.9703253e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001010001111110100111010011000;
		b = 32'b10111010010101110001100100001011;
		correct = 32'b11000101001000001011110110111001;
		#400 //3134374.0 * -0.0008205331 = -2571.8577
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110011111101101111001001000101;
		b = 32'b00010101000111100111100110100101;
		correct = 32'b11001001100110001101111011011110;
		#400 //-3.9130214e+31 * 3.2003807e-26 = -1252315.8
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000101110011101001111101101011;
		b = 32'b00001100000000001001010010011110;
		correct = 32'b10010010010011111000111101010010;
		#400 //-6611.9272 * 9.905484e-32 = -6.549434e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000111110001001101000101010101;
		b = 32'b00110001011101010100100111000001;
		correct = 32'b10111001101111001001010100001010;
		#400 //-100770.664 * 3.5694117e-09 = -0.00035969197
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001010111010000111111111011101;
		b = 32'b00100110001001010101000110011010;
		correct = 32'b10110001100101100010010010000110;
		#400 //-7618542.5 * 5.7356465e-16 = -4.369727e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001100111010101010111010101111;
		b = 32'b01010100001001000111100100101010;
		correct = 32'b10100001100101101100011011111011;
		#400 //-3.6158542e-31 * 2825629700000.0 = -1.0217065e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101100100100010101110101111100;
		b = 32'b01010101111100011101011001101101;
		correct = 32'b11000011000010010101001011000100;
		#400 //-4.1315267e-12 * 33237907000000.0 = -137.3233
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111110100101110011011010111101;
		b = 32'b10101110000100100110110100100100;
		correct = 32'b11101101001011001111101101011111;
		#400 //1.0049882e+38 * -3.3293493e-11 = -3.345957e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101101110111111100101110001111;
		b = 32'b00100000101001001000110111110011;
		correct = 32'b11001111000011111101101001111111;
		#400 //-8.6576556e+27 * 2.7876615e-19 = -2413461200.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011011101111000011001011000010;
		b = 32'b00011111101011111000001101101000;
		correct = 32'b10111100000000010000011101001101;
		#400 //-1.0594621e+17 * 7.4332776e-20 = -0.007875276
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101011000110110101110110110101;
		b = 32'b10001011101000110000111010110110;
		correct = 32'b10110111010001011110101100110000;
		#400 //1.8782602e+26 * -6.280745e-32 = -1.1796874e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110000111000111001101001101;
		b = 32'b01110000010010001010010000010001;
		correct = 32'b11100110111101010011110010110001;
		#400 //-2.3312925e-06 * 2.4838138e+29 = -5.7904967e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100011000011011001010100000010;
		b = 32'b01000011100101001100000101001000;
		correct = 32'b00100111001001001000101000010101;
		#400 //7.675179e-18 * 297.51 = 2.2834426e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111100000000001110000110111011;
		b = 32'b01101010100101100100100000111101;
		correct = 32'b11100111000101110101000101000100;
		#400 //-0.007866318 * 9.084e+25 = -7.145764e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101111110101000111100010000010;
		b = 32'b11001111000000000011111011010110;
		correct = 32'b11111111010101001110000011010000;
		#400 //1.3151301e+29 * -2151601700.0 = -2.8296363e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001001000100110100000101101100;
		b = 32'b10111011010011100101000011101001;
		correct = 32'b01000100111011010101101001011111;
		#400 //-603158.75 * -0.0031481332 = 1898.8241
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110100100110110100010011111110;
		b = 32'b01100001011011100000010011010100;
		correct = 32'b01010110100100000101110100010010;
		#400 //2.8921198e-07 * 2.7441706e+20 = 79364700000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010000111000101111011000110111;
		b = 32'b01111000000111101101110011001011;
		correct = 32'b11001001100011001101011110110110;
		#400 //-8.9520636e-29 * 1.2888455e+34 = -1153782.8
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100100011111110000001001011000;
		b = 32'b10100110011110110110100110011001;
		correct = 32'b01001011011110100111000001111101;
		#400 //-1.8816354e+22 * -8.722623e-16 = 16412797.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000010001100001000100100001010;
		b = 32'b00100110110101000011000100111111;
		correct = 32'b10101001100100100101001101110010;
		#400 //-44.133827 * 1.4723803e-15 = -6.498178e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100111110110000000111001110110;
		b = 32'b10100111101001100101011110101010;
		correct = 32'b00010000000011000110001101011101;
		#400 //-5.996772e-15 * -4.61693e-15 = 2.7686678e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111100000101111111010001100110;
		b = 32'b10101101011110001000010000001111;
		correct = 32'b10101010000100111000001100100110;
		#400 //0.009274578 * -1.4126491e-11 = -1.3101724e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000000110010010001111011001100;
		b = 32'b00111010001010001111011000111100;
		correct = 32'b00111011100001001011110110101001;
		#400 //6.2850094 * 0.0006445383 = 0.0040509296
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000011111010101100100010101111;
		b = 32'b11010111101000110110010111101000;
		correct = 32'b00011100000101011101101100111101;
		#400 //-1.3799359e-36 * -359316160000000.0 = 4.9583323e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000010010001010001110100010100;
		b = 32'b00110010110010100000101110000101;
		correct = 32'b00110101100110111001000111010000;
		#400 //49.278397 * 2.3521133e-08 = 1.1590837e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001000100100010100001110000101;
		b = 32'b01010001011010010110110101001010;
		correct = 32'b11011010100001000111010001111000;
		#400 //-297500.16 * 62660060000.0 = -1.8641378e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011100101111011100010110011101;
		b = 32'b11011011011111001101010100110010;
		correct = 32'b00111000101110110110110010010001;
		#400 //-1.2558053e-21 * -7.1166105e+16 = 8.937077e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100000101101011001010100101101;
		b = 32'b11010101001101110001111100100100;
		correct = 32'b11110110100000011110001110111010;
		#400 //1.0467531e+20 * -12584023000000.0 = -1.3172366e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010101100001111110010110111111;
		b = 32'b11011100011000100100100111110111;
		correct = 32'b00110010011100000100000000101101;
		#400 //-5.488854e-26 * -2.5477868e+17 = 1.39844305e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100100100110100011101010001110;
		b = 32'b10111010000001000000101011001100;
		correct = 32'b11011111000111110001100101100101;
		#400 //2.2760143e+22 * -0.0005037009 = -1.1464305e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100000110000110101101101111011;
		b = 32'b10011110001000011011011011111101;
		correct = 32'b00111111011101101101000001011001;
		#400 //-1.1261584e+20 * -8.56111e-21 = 0.96411663
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101000000110001110101001011110;
		b = 32'b01110000001111100111111001101010;
		correct = 32'b11011000111000111001001011101001;
		#400 //-8.488515e-15 * 2.358199e+29 = -2001760900000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011001000100111000001101000100;
		b = 32'b01000101101001001000101100101011;
		correct = 32'b11011111001111011010000010010001;
		#400 //-2595071900000000.0 * 5265.396 = -1.3664081e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110100000100111101110110101;
		b = 32'b01001100101011011011110011100001;
		correct = 32'b11000011101100010001101110111110;
		#400 //-3.8887033e-06 * 91088650.0 = -354.21674
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000001010101001000001111110111;
		b = 32'b11100101000100110011011010011101;
		correct = 32'b01100110111101000110101000111010;
		#400 //-13.282218 * -4.3449707e+22 = 5.7710848e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100010001001101001010001011101;
		b = 32'b11110110000110010000010001011100;
		correct = 32'b01011000110001110010001100000100;
		#400 //-2.2575738e-18 * -7.758885e+32 = 1751625600000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110000010101010110010001000110;
		b = 32'b10001000100001100001111001101111;
		correct = 32'b00111001010111111001011110110110;
		#400 //-2.6416612e+29 * -8.071987e-34 = 0.00021323454
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001010010100101011010011110001;
		b = 32'b00111101000111100111001011110110;
		correct = 32'b01001000000000100110101001001100;
		#400 //3452220.2 * 0.038683854 = 133545.19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101100100010111110001100001000;
		b = 32'b01010001101101101000101110101011;
		correct = 32'b11111110110001110111111101110011;
		#400 //-1.3529025e+27 * 98003410000.0 = -1.3258906e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010000010110100000110010111;
		b = 32'b10100001010100011001100111100101;
		correct = 32'b00011011111001000000100010000110;
		#400 //-0.0005312203 * -7.101563e-19 = 3.7724944e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000111011100110110110010011110;
		b = 32'b10111101011110010111100110111111;
		correct = 32'b10000101011011010011100001101010;
		#400 //1.8313208e-34 * -0.06090712 = -1.1154048e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010101000110001010000001101010;
		b = 32'b01001101100011110001110011101010;
		correct = 32'b00100011001010101010010110110001;
		#400 //3.08227e-26 * 300129600.0 = 9.250805e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010000111010010001000110011110;
		b = 32'b10111001111110111011100111101101;
		correct = 32'b00001011011001010010110110001011;
		#400 //-9.192944e-29 * -0.00048012976 = 4.4138058e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000000010101000010100101001100;
		b = 32'b11011001100001010000011110110100;
		correct = 32'b10011010001011101110111111110011;
		#400 //7.728996e-39 * -4680580000000000.0 = -3.6176186e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010000010101110001110101100111;
		b = 32'b10010100111101010001000001100010;
		correct = 32'b00100101110011011110110011101000;
		#400 //-14436113000.0 * -2.474514e-26 = 3.5722365e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010110100101001010011101101011;
		b = 32'b11001110111010001001010110011100;
		correct = 32'b01100110000001110000111010011001;
		#400 //-81723390000000.0 * -1951059500.0 = 1.5944719e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000011101011111100111101001011;
		b = 32'b01000000011101111101101000111000;
		correct = 32'b11000100101010100011011011011110;
		#400 //-351.61948 * 3.872694 = -1361.7146
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100000110100101010001110000;
		b = 32'b00100110001010001010001100110101;
		correct = 32'b00101010110010110101001110011010;
		#400 //617.31934 * 5.8507896e-16 = 3.6118054e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110011011001111111111000001010;
		b = 32'b11111001001010000111101101101101;
		correct = 32'b01101101000110001010111010010000;
		#400 //-5.4014926e-08 * -5.467558e+34 = 2.9532972e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001011110011101101101000110111;
		b = 32'b01000011110010100110101100111111;
		correct = 32'b10010000001000111000111011011000;
		#400 //-7.9676647e-32 * 404.83786 = -3.2256125e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000000100101001001110101011100;
		b = 32'b00001011001111011001110111000100;
		correct = 32'b10001100010111000010011110000110;
		#400 //-4.644209 * 3.6518766e-32 = -1.6960077e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000000101011110011101101011100;
		b = 32'b00010001110001001111010001101100;
		correct = 32'b00010011000001101101000011000001;
		#400 //5.475996 * 3.1073984e-28 = 1.7016101e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011100000101110111000010000110;
		b = 32'b10101010000010000010010010110001;
		correct = 32'b11000110101000010001001011110111;
		#400 //1.7050577e+17 * -1.2091956e-13 = -20617.482
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110010010100001010100011101000;
		b = 32'b10011111001010110101101011110111;
		correct = 32'b00010010000010111010101011111000;
		#400 //-1.2145598e-08 * -3.6285903e-20 = 4.40714e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111001000110110000001010111101;
		b = 32'b11000011000110010101011000011011;
		correct = 32'b01111100101110011011000110001100;
		#400 //-5.0303847e+34 * -153.33635 = 7.713408e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100111111100000111010110010101;
		b = 32'b00111110010101001110001101101001;
		correct = 32'b00100110110001111111011011111010;
		#400 //6.6740864e-15 * 0.20789875 = 1.3875342e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110101110011001010001000010001;
		b = 32'b10100010101011011010101101000001;
		correct = 32'b10011001000010101101001001101010;
		#400 //1.5246352e-06 * -4.7073066e-18 = -7.1769256e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101100100000110111010110001101;
		b = 32'b00101000101011001110010110101110;
		correct = 32'b11010101101100011001000111011000;
		#400 //-1.2713952e+27 * 1.9195444e-14 = -24404994000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000101010110110000001011000001;
		b = 32'b10100101000101110010000111111101;
		correct = 32'b10101011000000010100101110110100;
		#400 //3504.172 * -1.3108678e-16 = -4.5935066e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001001011111101011000111110000;
		b = 32'b00101010101110001111110001010111;
		correct = 32'b10110100101110000000101011110010;
		#400 //-1043231.0 * 3.2860062e-13 = -3.4280635e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001010100111111110110001000101;
		b = 32'b01110010100000111000011001110011;
		correct = 32'b01111101101001000101001111001010;
		#400 //5240354.5 * 5.2102497e+30 = 2.7303556e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010011110011010110011011101001;
		b = 32'b11000100110100101000000100100111;
		correct = 32'b11011001001010001110011000001011;
		#400 //1764389700000.0 * -1684.036 = -2971295700000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010100100101101110100000011100;
		b = 32'b01001101001101010010101000000100;
		correct = 32'b01100010010101011001010111000000;
		#400 //5185114000000.0 * 189964350.0 = 9.849868e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110111011010110000110000111110;
		b = 32'b10001101111000010011010111110011;
		correct = 32'b01000101110011101100011101001011;
		#400 //-4.7673362e+33 * -1.3879683e-30 = 6616.9116
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000110101001110001000110100101;
		b = 32'b01010001001100110100001101000111;
		correct = 32'b00011000011010011111101001111101;
		#400 //6.2844344e-35 * 48120490000.0 = 3.0241008e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000010001100001100101111010;
		b = 32'b11000111100011010111001101010000;
		correct = 32'b00111000010110101110101010000111;
		#400 //-7.2068185e-10 * -72422.625 = 5.219367e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001000110001101110000101100001;
		b = 32'b11101101101111000111101011010111;
		correct = 32'b11110111000100100110110011110010;
		#400 //407307.03 * -7.291461e+27 = -2.9698633e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011011110001100111101001100001;
		b = 32'b00010111110110101101011110001001;
		correct = 32'b10110100001010011010101101010010;
		#400 //-1.11733205e+17 * 1.4142329e-24 = -1.5801677e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011101111000100100101100100110;
		b = 32'b11011110101000000111101001101100;
		correct = 32'b00111101000011011101101100101111;
		#400 //-5.9899404e-21 * -5.781837e+18 = 0.034632858
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110111010111001100001100110000;
		b = 32'b00011110001100101110101101101111;
		correct = 32'b00010110000110100100101010111110;
		#400 //1.31584675e-05 * 9.471928e-21 = 1.2463605e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111100011111111000001100001001;
		b = 32'b10011110001100100100001110000010;
		correct = 32'b01011011001100011110110001111101;
		#400 //-5.3067736e+36 * -9.437202e-21 = 5.0081092e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110000011011101011100011010;
		b = 32'b10111001110000110111100011111110;
		correct = 32'b00110000010110001001101111000101;
		#400 //-2.1135843e-06 * -0.00037283445 = 7.8801704e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111001010101100010111111010111;
		b = 32'b10110110010000111011100100101110;
		correct = 32'b01110000001000111100000101100000;
		#400 //-6.9507615e+34 * -2.9165053e-06 = 2.0271933e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000000110001100001100110000100;
		b = 32'b11011101001000101111011111000010;
		correct = 32'b11011110011111000011011110111101;
		#400 //6.1906147 * -7.3394174e+17 = -4.5435507e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110000100000011101101001010010;
		b = 32'b10001000011000001110001101110000;
		correct = 32'b10111001011001000010010011001010;
		#400 //3.215e+29 * -6.76749e-34 = -0.0002175748
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011101000010110010110100111011;
		b = 32'b01100101100101000010000110011001;
		correct = 32'b01000011001000010001000011010100;
		#400 //1.841988e-21 * 8.744125e+22 = 161.06573
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000101101111101011101110010;
		b = 32'b10111100110001110111010000110110;
		correct = 32'b00101110000011110011101111101110;
		#400 //-1.3376236e-09 * -0.024347406 = 3.2567664e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000110101100110010111101010101;
		b = 32'b11110101101101010100101100001111;
		correct = 32'b11111100111111011100101000000001;
		#400 //22935.666 * -4.5963286e+32 = -1.0541986e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011111110001101010110110101;
		b = 32'b11010000111001010100010100100101;
		correct = 32'b01011101010111101101101001100000;
		#400 //-32615274.0 * -30772111000.0 = 1.0036408e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010001001110001010100001110111;
		b = 32'b01000100111000000000111001111011;
		correct = 32'b00010110101000011001110111011010;
		#400 //1.4566953e-28 * 1792.4525 = 2.611057e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111010011001101001000000011111;
		b = 32'b01110000110100100001001001110110;
		correct = 32'b01101011101111010011001011011010;
		#400 //0.00087952794 * 5.2011336e+29 = 4.5745424e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010001101001110001100101000101;
		b = 32'b10101110011101011111010111000011;
		correct = 32'b10000000101000001000101110011010;
		#400 //2.6363528e-28 * -5.592483e-11 = -1.4743759e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001000011110100110001010011010;
		b = 32'b11000011010001100000010010010111;
		correct = 32'b00001100010000011010110011000000;
		#400 //-7.5347544e-34 * -198.01793 = 1.4920164e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001010001100100100111011111100;
		b = 32'b10110110011100010100011111001001;
		correct = 32'b00000001001010000000111001011011;
		#400 //-8.5852436e-33 * -3.5953583e-06 = 3.0867026e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011100001101000000111101000101;
		b = 32'b01001000010110010110110110001100;
		correct = 32'b11100101000110001110110111111110;
		#400 //-2.0272914e+17 * 222646.19 = -4.513687e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111010111010110001101001011101;
		b = 32'b00100010010101101011000000101111;
		correct = 32'b11011101110001010010100111010111;
		#400 //-6.1036224e+35 * 2.9095679e-18 = -1.7758904e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100001010011101100011001111101;
		b = 32'b00100000111100110101001000011000;
		correct = 32'b01000010110001001000100010111000;
		#400 //2.3839574e+20 * 4.1220126e-19 = 98.26703
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110110111101101001000010100101;
		b = 32'b11101000100000111000001110111001;
		correct = 32'b11011111111111010101010111000101;
		#400 //7.34821e-06 * -4.968479e+24 = -3.6509427e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110000101001111111010100100101;
		b = 32'b01101001010101000000001001100101;
		correct = 32'b01011010100010110001100010010101;
		#400 //1.2220523e-09 * 1.6018974e+25 = 1.9576025e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100110111111011000110111010001;
		b = 32'b10011101010100100001110101111011;
		correct = 32'b10000100110100000001101110001000;
		#400 //1.7593841e-15 * -2.780851e-21 = -4.892585e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010111001101101000011001010111;
		b = 32'b01011010001000011010101001101000;
		correct = 32'b10110001111001101000011111111000;
		#400 //-5.897693e-25 * 1.1376209e+16 = -6.709339e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010010011001111010010000111111;
		b = 32'b01101100101101101010110111011110;
		correct = 32'b00111111101001010100110000011000;
		#400 //7.3093197e-28 * 1.7667645e+27 = 1.2913847
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110001000010001010100100101001;
		b = 32'b10010001010000001101100000011100;
		correct = 32'b01000010110011011110010001111001;
		#400 //-6.767114e+29 * -1.5212723e-28 = 102.946236
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101110101011111011101001010000;
		b = 32'b00010111000011100100110001000000;
		correct = 32'b11000110010000110101101101011111;
		#400 //-2.7192557e+28 * 4.5978916e-25 = -12502.843
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000011111001111110101000010010;
		b = 32'b11010100011111110111011001010001;
		correct = 32'b10011000111001110110110101010111;
		#400 //1.36307e-36 * -4388806700000.0 = -5.9822505e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101101001101010110101000100010;
		b = 32'b11110010101011001000101011010100;
		correct = 32'b01100000011101001000101101100001;
		#400 //-1.0312225e-11 * -6.8351046e+30 = 7.048514e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101101101010001101011000110000;
		b = 32'b10001110000100010001011101110011;
		correct = 32'b10111100001111110110000110010001;
		#400 //6.5315523e+27 * -1.788392e-30 = -0.0116809765
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011000111100000110011100010110;
		b = 32'b11011010000010100101110110100100;
		correct = 32'b01110011100000011110111110000001;
		#400 //-2114604300000000.0 * -9736626000000000.0 = 2.0589112e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011100010000101001101011111001;
		b = 32'b11010110111101000100000101010100;
		correct = 32'b01110011101110011010110101011111;
		#400 //-2.1910616e+17 * -134280710000000.0 = 2.9421732e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100000111011000110110011011110;
		b = 32'b00111110100101110100010100111011;
		correct = 32'b00100000000010111011010000100111;
		#400 //4.0051997e-19 * 0.29545006 = 1.1833365e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100000111000000111000100111101;
		b = 32'b11001100010111001110110001010010;
		correct = 32'b11101101110000011011000010000001;
		#400 //1.293822e+20 * -57913670.0 = -7.4929984e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000101000000100101111011111100;
		b = 32'b11011111100011001110011100011101;
		correct = 32'b01100101000011111000001101001001;
		#400 //-2085.9365 * -2.0306232e+19 = 4.235751e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101100011010001001000001001001;
		b = 32'b10000101000001001010100100001000;
		correct = 32'b10110001111100010000011111101000;
		#400 //1.1246086e+27 * -6.237656e-36 = -7.014922e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101010111101001110010001000100;
		b = 32'b00010000001101001111100101110010;
		correct = 32'b00111011101011010001111100011111;
		#400 //1.4802793e+26 * 3.5690906e-29 = 0.005283251
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011110010101111101000010110111;
		b = 32'b11001110001111000000111100001010;
		correct = 32'b00101101000111101000100111110100;
		#400 //-1.14251664e-20 * -788775550.0 = 9.011892e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000011010001100001000110010000;
		b = 32'b01111101100101111010011010111010;
		correct = 32'b01000001011010101010101010110110;
		#400 //5.820713e-37 * 2.519739e+37 = 14.666677
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111011111101011000000010100000;
		b = 32'b10001100011110010000001110100001;
		correct = 32'b10001000111011101100110110010111;
		#400 //0.00749214 * -1.9183354e-31 = -1.4372438e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101111010100001010100100101010;
		b = 32'b00011011001010101010010000000010;
		correct = 32'b10001011000010110001011000000100;
		#400 //-1.8977589e-10 * 1.4115064e-22 = -2.678699e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001100000111110001000010010001;
		b = 32'b11110101111100111110101110001010;
		correct = 32'b01000010100101111000111100010100;
		#400 //-1.22539e-31 * -6.1841086e+32 = 75.77945
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100001001101011011111110000110;
		b = 32'b00111000000111000010001101000011;
		correct = 32'b00011001110111011011001101111101;
		#400 //6.1578665e-19 * 3.722614e-05 = 2.2923359e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110101001010010111111000000001;
		b = 32'b10101001000111110101110000100011;
		correct = 32'b10011110110100110000010010000110;
		#400 //6.3140766e-07 * -3.5385008e-14 = -2.2342365e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111010001111100010010111110101;
		b = 32'b01011011010001111101000011111000;
		correct = 32'b01010110000101000110101010111000;
		#400 //0.0007253581 * 5.6243284e+16 = 40796520000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100001010101011001001111110000;
		b = 32'b01000011011011011000111100010011;
		correct = 32'b10100101010001100011000101010011;
		#400 //-7.2363e-19 * 237.55888 = -1.7190474e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010010010000101110100001101000;
		b = 32'b11010100111011101111011000100010;
		correct = 32'b01100111101101011110111101110110;
		#400 //-209280700000.0 * -8210653000000.0 = 1.7183312e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011010011100010000100011010011;
		b = 32'b11010110011011110111010011010100;
		correct = 32'b10110001011000010111010100111101;
		#400 //4.984476e-23 * -65821263000000.0 = -3.2808452e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000001110110111111001011111001;
		b = 32'b10100100101111101011000101011111;
		correct = 32'b10100111001000111101011010111001;
		#400 //27.493639 * -8.2699843e-17 = -2.2737196e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001100111100100101011110011100;
		b = 32'b10100100110011000111111100111011;
		correct = 32'b00110010010000011001011001000010;
		#400 //-127057120.0 * -8.8686434e-17 = 1.1268243e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001001101111010010101000111000;
		b = 32'b10111110000101101101101000110100;
		correct = 32'b11001000010111101110111111110010;
		#400 //1549639.0 * -0.14731675 = -228287.78
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010110000011100111011111001000;
		b = 32'b01111000101001010001010101111011;
		correct = 32'b11001111001101111011111001010000;
		#400 //-1.1508465e-25 * 2.6786396e+34 = -3082702800.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101000100101010011100100110011;
		b = 32'b11001101000110000110110011100001;
		correct = 32'b01110110001100011011001011011011;
		#400 //-5.637502e+24 * -159829520.0 = 9.010392e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101010111110000111100001110001;
		b = 32'b00010101101110011110011110100110;
		correct = 32'b11000001001101000110111111011111;
		#400 //-1.5019119e+26 * 7.508638e-26 = -11.277312
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011010100000100111001000101000;
		b = 32'b10100000011001000001000101101100;
		correct = 32'b00111011011010000110110100011000;
		#400 //-1.8358632e+16 * -1.9318116e-19 = 0.0035465416
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111001000100010101100011010111;
		b = 32'b10011110100001111111111001100001;
		correct = 32'b01011000000110100110110010001101;
		#400 //-4.716781e+34 * -1.439889e-20 = 679164050000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010010000111011011010110001111;
		b = 32'b01100100010110010011001010101011;
		correct = 32'b01110111000001011100111000011101;
		#400 //169338980000.0 * 1.6026378e+22 = 2.7138905e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101000010110011100101000101000;
		b = 32'b00000010101010110101101000011101;
		correct = 32'b10101011100100011100011010110010;
		#400 //-4.1139306e+24 * 2.5177914e-37 = -1.0358019e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011000110001110101011110011010;
		b = 32'b11110001001101111111101110100001;
		correct = 32'b01001010100011110100001110001111;
		#400 //-5.152875e-24 * -9.110393e+29 = 4694471.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110011110101011010100101101110;
		b = 32'b01110010000111010101101110111111;
		correct = 32'b01100110100000110101010101111011;
		#400 //9.9494045e-08 * 3.116804e+30 = 3.1010342e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011100110110111101000010101101;
		b = 32'b00010111010001111101001000111100;
		correct = 32'b10110100101010111001001110111011;
		#400 //-4.949797e+17 * 6.456572e-25 = -3.195872e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011000110011011001001001101111;
		b = 32'b10111111011100011010011001011011;
		correct = 32'b10011000110000100000110001110001;
		#400 //5.313912e-24 * -0.94394463 = -5.0160387e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001000100011111010110110000101;
		b = 32'b01001000101010001111110011000100;
		correct = 32'b10010001101111011010111101111000;
		#400 //-8.647294e-34 * 346086.12 = -2.9927083e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110101010000001001101101101010;
		b = 32'b10110001000110111010100011010111;
		correct = 32'b11100110111010100011101001000010;
		#400 //2.4415849e+32 * -2.2651443e-09 = -5.530542e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110100100100000110101111111010;
		b = 32'b10010100100011000101011111111010;
		correct = 32'b00001001100111100101100101011101;
		#400 //-2.6900653e-07 * -1.4171088e-26 = 3.8121153e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010001100100100111011101100101;
		b = 32'b00111101101001100110011010011010;
		correct = 32'b01001111101111100110100000111110;
		#400 //78633540000.0 * 0.081250384 = 6389005300.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101100011010101000100000001110;
		b = 32'b00111011001000001011011101001100;
		correct = 32'b11101000000100110011110011110110;
		#400 //-1.1341246e+27 * 0.0024523316 = -2.7812496e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111100011001000101011000101010;
		b = 32'b00100001111110000111100100110001;
		correct = 32'b11011110110111011001111110010001;
		#400 //-4.7423652e+36 * 1.6837213e-18 = -7.984821e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010010110101101001011111001000;
		b = 32'b01010001001110011111111100101100;
		correct = 32'b01100100100110111110100110010110;
		#400 //460834730000.0 * 49928126000.0 = 2.3008616e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110010111000010010001010001101;
		b = 32'b11000100111110110001011011000100;
		correct = 32'b00111000010111001101000011100110;
		#400 //-2.620916e-08 * -2008.7114 = 5.264664e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000001000100111100000001011011;
		b = 32'b01100011001011110010010011110101;
		correct = 32'b00100100110010100010101110100101;
		#400 //2.7137644e-38 * 3.2308432e+21 = 8.767747e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000000000010100101110111111001;
		b = 32'b01010011010110001110011100000001;
		correct = 32'b00010010100011001000101001001111;
		#400 //9.52066e-40 * 931588540000.0 = 8.869338e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100000101110101110101000001101;
		b = 32'b01110011000010011011101000001111;
		correct = 32'b01010100010010010001111000110100;
		#400 //3.1664507e-19 * 1.0911841e+31 = 3455180600000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001011010111100011101110101000;
		b = 32'b11011111000111011000101000110101;
		correct = 32'b10101011000010001100001010010000;
		#400 //4.2800525e-32 * -1.1351944e+19 = -4.8586916e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011010011111110111000011110110;
		b = 32'b10110101010101011110000111001111;
		correct = 32'b10010000010101010110101001001110;
		#400 //5.2824013e-23 * -7.967728e-07 = -4.2088737e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001010101001110011100000111101;
		b = 32'b10001011001001010100100110000000;
		correct = 32'b10010110010101111110111010000100;
		#400 //5479454.5 * -3.183314e-32 = -1.7442824e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101101000100101010111011111010;
		b = 32'b00000110101110001111111100001100;
		correct = 32'b10110100010100111111111111001110;
		#400 //-2.8372716e+27 * 6.9587865e-35 = -1.9743968e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000011100111111110111001111101;
		b = 32'b01010000001101001001000011111000;
		correct = 32'b10010100011000011001110010000010;
		#400 //-9.399934e-37 * 12117598000.0 = -1.1390463e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000101101100111000101110110010;
		b = 32'b11101100110011011000000010110011;
		correct = 32'b10110011000100000010000100100001;
		#400 //1.6884395e-35 * -1.9875005e+27 = -3.3557743e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100101010100010100100111101001;
		b = 32'b10101000010110001010111111011010;
		correct = 32'b00001110001100010010011000100000;
		#400 //-1.8152902e-16 * -1.202854e-14 = 2.183529e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011010000100101001101000110010;
		b = 32'b11000101100000011001110000111010;
		correct = 32'b11100000000101000111001001010101;
		#400 //1.0316222e+16 * -4147.5283 = -4.278682e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010001101101001110110000101010;
		b = 32'b01100011110010011110100101100000;
		correct = 32'b01110110000011101011001001011100;
		#400 //97132040000.0 * 7.449224e+21 = 7.235583e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110101111110110000111010011;
		b = 32'b11011101110001010011001011011111;
		correct = 32'b01010101000100110110110001001111;
		#400 //-5.703632e-06 * -1.7762081e+18 = 10130837000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111110010010101110001000101000;
		b = 32'b10010101101011011001011001001100;
		correct = 32'b11010100100010011001000111110010;
		#400 //6.741958e+37 * -7.011127e-26 = -4726872600000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111000101010001000011110010000;
		b = 32'b10000101110010011101100111101011;
		correct = 32'b10111111000001001110000111100110;
		#400 //2.7345481e+34 * -1.8982e-35 = -0.51907194
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111111110110110111101011011100;
		b = 32'b01111001010111100000101101001111;
		correct = 32'b11111001101111100101111000111101;
		#400 //-1.7146869 * 7.2057454e+34 = -1.2355597e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000110111110100011011011010111;
		b = 32'b11100100000111111010100011000100;
		correct = 32'b01101011100111000000110100000011;
		#400 //-32027.42 * -1.1780773e+22 = 3.7730775e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101001100001101110111111010101;
		b = 32'b11001101011101001000110010011100;
		correct = 32'b00110111100000001110011010110100;
		#400 //-5.9923996e-14 * -256428480.0 = 1.5366219e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000000000011111111111111100110;
		b = 32'b10100001110001101010011100110100;
		correct = 32'b00100010010111110111101111110010;
		#400 //-2.2499938 * -1.346126e-18 = 3.0287752e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010101010110010000111000101111;
		b = 32'b10110001001001011000110101101100;
		correct = 32'b10000111000011000101111000001101;
		#400 //4.383399e-26 * -2.409105e-09 = -1.0560068e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100011011101100000100001010010;
		b = 32'b11001101000011001010101010111001;
		correct = 32'b10110001000001110011000010100000;
		#400 //1.3337449e-17 * -147499920.0 = -1.9672726e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111110000110000100110110110000;
		b = 32'b10110110001100100010110011110111;
		correct = 32'b01110100110101000000000110001001;
		#400 //-5.061151e+37 * -2.655024e-06 = 1.3437476e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010100011111011101010101100001;
		b = 32'b10111110111000000110100110011000;
		correct = 32'b10010011110111101000001101101000;
		#400 //1.2815317e-26 * -0.43830562 = -5.6170255e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000010001101011000011000110001;
		b = 32'b11100010101111100000111001001101;
		correct = 32'b11100101100001101100001110111100;
		#400 //45.381046 * -1.7529559e+21 = -7.955097e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011001010000001000100111010110;
		b = 32'b10001111100100110110100001010011;
		correct = 32'b00101001010111011011101100111001;
		#400 //-3387171700000000.0 * -1.4535503e-29 = 4.9234247e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111101111111100110011011000011;
		b = 32'b10000110000001101111000001011110;
		correct = 32'b01000100100001100001100010101000;
		#400 //-4.2269685e+37 * -2.5379193e-35 = 1072.7705
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000001001110010001111111010101;
		b = 32'b01001100011001010111010100001110;
		correct = 32'b00001110001001011110111000011111;
		#400 //3.4001972e-38 * 60150840.0 = 2.0452471e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100010010010111000111110010111;
		b = 32'b01111110101001011101011110011001;
		correct = 32'b11100001100000111101111011111100;
		#400 //-2.7587646e-18 * 1.1022103e+38 = -3.040739e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000001101110001111101100110001;
		b = 32'b10110101011000100100000011111101;
		correct = 32'b10110111101000110111110010110111;
		#400 //23.122652 * -8.428613e-07 = -1.9489189e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011110101100110110101010011100;
		b = 32'b00000001000010000000001011010100;
		correct = 32'b00100000001111101010010100111101;
		#400 //6.4641586e+18 * 2.4981284e-38 = 1.6148299e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011101010010000001110100011101;
		b = 32'b01100110111000011011010101100000;
		correct = 32'b11000100101100000110111101011110;
		#400 //-2.648483e-21 * 5.3293912e+23 = -1411.4802
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010110101011011001111111110111;
		b = 32'b01110010010111000001011110010000;
		correct = 32'b01001001100101010100010101110011;
		#400 //2.805061e-25 * 4.359372e+30 = 1222830.4
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110000000101000010110001010101;
		b = 32'b10001111000101011011101000111101;
		correct = 32'b10111111101011010101001100110010;
		#400 //1.834295e+29 * -7.382135e-30 = -1.3541014
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101111001100011101111011111110;
		b = 32'b10010100000010010000011111001001;
		correct = 32'b10000011101111100110101101111101;
		#400 //1.6177279e-10 * -6.918268e-27 = -1.1191874e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000101110110111010111111001101;
		b = 32'b11001010111010110001011100011001;
		correct = 32'b11010001010010011011111000110011;
		#400 //7029.975 * -7703436.5 = -54154965000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011000000011100111101010001111;
		b = 32'b10101010010001111111101001001001;
		correct = 32'b01000010110111101001100100100011;
		#400 //-626628150000000.0 * -1.7761586e-13 = 111.299095
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000010101000110001101011011001;
		b = 32'b01111001011100111011110101101111;
		correct = 32'b11111100100110110100101100101110;
		#400 //-81.55244 * 7.9098144e+34 = -6.450647e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010101100100110011001110110110;
		b = 32'b11111110000001110100010001001010;
		correct = 32'b01010100000110111000111100010011;
		#400 //-5.945441e-26 * -4.495009e+37 = 2672481300000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100011001110001011000010011111;
		b = 32'b00111111001000000011000001101111;
		correct = 32'b10100010111001110010001010101001;
		#400 //-1.0012061e-17 * 0.62573904 = -6.2649373e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100011001100101101011101111011;
		b = 32'b01110001000111110001100001110100;
		correct = 32'b11010100110111100100100111010101;
		#400 //-9.695029e-18 * 7.8780286e+29 = -7637771500000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000000100101100010100110010110;
		b = 32'b00111100011111000001100100010011;
		correct = 32'b10111101100100111101111110100101;
		#400 //-4.6925764 * 0.015386838 = -0.07220391
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111111000101100010101011110100;
		b = 32'b11101100100010100000100100010101;
		correct = 32'b11101100001000011111000011110111;
		#400 //0.5865929 * -1.3349972e+27 = -7.830999e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001000100101100011110000000111;
		b = 32'b01110011011100110111101101000000;
		correct = 32'b01111100100011101110001101001111;
		#400 //307680.22 * 1.9290588e+31 = 5.935332e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001111110110001001111011100011;
		b = 32'b01000000111011000101111110001011;
		correct = 32'b00010001010010000000001101010010;
		#400 //2.1360445e-29 * 7.386663 = 1.5778241e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110110101101011111011110010011;
		b = 32'b11011110001100000110111110111001;
		correct = 32'b11010101011110101101001100111110;
		#400 //5.423042e-06 * -3.178396e+18 = -17236574000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101001101001101100101111011000;
		b = 32'b01101101110010000111000010000111;
		correct = 32'b01011000000000101001100010010010;
		#400 //7.407242e-14 * 7.75413e+27 = 574367200000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111100000100010011001111010011;
		b = 32'b00100100101011011110010111111010;
		correct = 32'b00100001010001010100010011101101;
		#400 //0.0088624535 * 7.5416386e-17 = 6.683742e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101101010100110111001111010101;
		b = 32'b00100100101001110111000000001111;
		correct = 32'b11010010100010100100110100011111;
		#400 //-4.0900856e+27 * 7.261454e-17 = -296999680000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010100011001001001001011100100;
		b = 32'b00110100001010001110100000000000;
		correct = 32'b01001001000101101100111110001011;
		#400 //3926867800000.0 * 1.573062e-07 = 617720.7
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100000111000100010110100010010;
		b = 32'b10110110011100000100011010101010;
		correct = 32'b00010111110101000100100010101111;
		#400 //-3.8315714e-19 * -3.5803919e-06 = 1.3718527e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001000011011101101011010001011;
		b = 32'b10000111110000000001100011110100;
		correct = 32'b00010000101100110011100000110000;
		#400 //-244570.17 * -2.8903615e-34 = 7.068962e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010101100101100111010010011001;
		b = 32'b01000011100110101001100001011001;
		correct = 32'b10011001101101011011011101011011;
		#400 //-6.0768476e-26 * 309.19022 = -1.8789018e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011001001000100001010010110011;
		b = 32'b01110111000110000011001111001101;
		correct = 32'b01010000110000001011101000101100;
		#400 //8.379384e-24 * 3.0870303e+33 = 25867411000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100111110011111111001011100111;
		b = 32'b00110100011111110100010110011101;
		correct = 32'b01011100110011110101101110000000;
		#400 //1.9640212e+24 * 2.3774051e-07 = 4.669274e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010110010110010001010001101000;
		b = 32'b10111100011101110110010110011001;
		correct = 32'b10010011010100011100100011010111;
		#400 //1.753556e-25 * -0.015099906 = -2.647853e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011100100011000111111011101000;
		b = 32'b00100110001101011010010001011010;
		correct = 32'b10000011010001110101111111011001;
		#400 //-9.297227e-22 * 6.301973e-16 = -5.859087e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010011110011011100001011100011;
		b = 32'b00100110100110101000000001001000;
		correct = 32'b10111010111110000101110010110000;
		#400 //-1767475900000.0 * 1.0720667e-15 = -0.0018948521
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010011110011101101100110000010;
		b = 32'b11010101001101011100011111000011;
		correct = 32'b10101001100100101110000100110010;
		#400 //5.221619e-27 * -12491848000000.0 = -6.5227676e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110011101101101010000000100100;
		b = 32'b00011111001010101011011000001011;
		correct = 32'b10010011011100111001000001101011;
		#400 //-8.504165e-08 * 3.6149483e-20 = -3.0742116e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011011110110110110010100011010;
		b = 32'b11100010001111001101010110001110;
		correct = 32'b00111110101000011101010101000100;
		#400 //-3.6295846e-22 * -8.70844e+20 = 0.3160802
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111101111110100010110101001000;
		b = 32'b00111111101011011111110111010001;
		correct = 32'b00111110001010100000100010100101;
		#400 //0.12215668 * 1.3593084 = 0.1660486
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001001101000110101000010111000;
		b = 32'b10001111110111101100100100111100;
		correct = 32'b00011010000011100010000001100000;
		#400 //-1337879.0 * -2.1968403e-29 = 2.9391064e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000011000110110101100110101101;
		b = 32'b11001001010011111100010111000111;
		correct = 32'b01001100111111000010101100001111;
		#400 //-155.3503 * -851036.44 = 132208760.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110001111001111000000000110111;
		b = 32'b10000010100001111011110000010101;
		correct = 32'b00110100111101010111110101100100;
		#400 //-2.2926733e+30 * -1.994442e-37 = 4.572604e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010001011101101011000111000011;
		b = 32'b10111110100001001001110110110111;
		correct = 32'b10010000011111111001011101001000;
		#400 //1.9460755e-28 * -0.25901577 = -5.0406426e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001001111101110100100110000010;
		b = 32'b00100100000000011101010011001110;
		correct = 32'b10101110011110101101001100110101;
		#400 //-2025776.2 * 2.815267e-17 = -5.703101e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001000111110111111010111110001;
		b = 32'b11011100001010001000111101101100;
		correct = 32'b00100101101001011110011010001111;
		#400 //-1.5164334e-33 * -1.8978196e+17 = 2.877917e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011101101000011100011110010000;
		b = 32'b10100010101101100101111000111011;
		correct = 32'b10000000111001100111111011011010;
		#400 //4.2822688e-21 * -4.943097e-18 = -2.116767e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011111111010100000101010111011;
		b = 32'b11011100010101111001001011100101;
		correct = 32'b01111100110001010001010101001111;
		#400 //-3.3728995e+19 * -2.4271453e+17 = 8.1865174e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011110100010000010101101101010;
		b = 32'b01100001011101011100100001001101;
		correct = 32'b01000000100000101011110000010111;
		#400 //1.4417516e-20 * 2.8336784e+20 = 4.08546
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000000110010001000000001010100;
		b = 32'b00100010001110001111101000010010;
		correct = 32'b10100011100100001110000000011000;
		#400 //-6.265665 * 2.5069036e-18 = -1.5707419e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011111011011101011010001001111;
		b = 32'b10000010110000000110001101100101;
		correct = 32'b10100010101100110110001111101001;
		#400 //1.720046e+19 * -2.8268914e-37 = -4.862383e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100110111111100111110010001001;
		b = 32'b10110101111001101010110001010111;
		correct = 32'b10011101011001010100111100110101;
		#400 //1.7658546e-15 * -1.7186493e-06 = -3.0348847e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001000100011111010000001010000;
		b = 32'b00011110101001000010010000011011;
		correct = 32'b10100111101110000010110111101010;
		#400 //-294146.5 * 1.7379108e-20 = -5.112004e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100111100110101011111100110111;
		b = 32'b00011111101011111110000000110100;
		correct = 32'b10000111110101001010000001111011;
		#400 //-4.29509e-15 * 7.4486296e-20 = -3.1992537e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011010111111101100101100110000;
		b = 32'b11101101001110101101111011100001;
		correct = 32'b11001000101110011111110101110101;
		#400 //1.05380205e-22 * -3.6146035e+27 = -380907.66
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101011000100011010100100111100;
		b = 32'b01110101011000110011110100000111;
		correct = 32'b11100001000000010100101111001010;
		#400 //-5.174921e-13 * 2.8805888e+32 = -1.490682e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010101101111111101001010100101;
		b = 32'b00010101100000110000110101011111;
		correct = 32'b10101011110001000110010110011111;
		#400 //-26363930000000.0 * 5.2931575e-26 = -1.3954843e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101011001001001110101110011010;
		b = 32'b10010100111111110111111101000000;
		correct = 32'b01000000101001001001100010101001;
		#400 //-1.9937643e+26 * -2.5798611e-26 = 5.1436353
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011100110111110111111000000110;
		b = 32'b11100000010001001111010011010101;
		correct = 32'b01111101101010111111001000111011;
		#400 //-5.0325987e+17 * -5.676881e+19 = 2.8569465e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101111111110010100111000000101;
		b = 32'b00000111001000111001000011100001;
		correct = 32'b10110111100111110100100111000100;
		#400 //-1.5431217e+29 * 1.2305333e-34 = -1.8988627e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011111000100111010110010111001;
		b = 32'b01001001100111101001000100110110;
		correct = 32'b00101001001101101111000010111100;
		#400 //3.1271334e-20 * 1298982.8 = 4.0620922e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111110011001001001101110111;
		b = 32'b00111111010111001011011011000000;
		correct = 32'b01000111101100000110000011000101;
		#400 //104742.93 * 0.86216354 = 90305.54
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100000111111110001100000111101;
		b = 32'b01001100111001100010101100101100;
		correct = 32'b11101110011001010101101011001100;
		#400 //-1.4705207e+20 * 120674660.0 = -1.7745458e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010010011001101111001100001011;
		b = 32'b00100000100111011100111111011100;
		correct = 32'b00110011100011100101111010010011;
		#400 //247980020000.0 * 2.6734384e-19 = 6.629593e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101110101001000000101001110001;
		b = 32'b01110101110100111000001110101100;
		correct = 32'b11100101000001111000100011111011;
		#400 //-7.459711e-11 * 5.3625257e+32 = -4.0002895e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111010000110000101101101011000;
		b = 32'b11000001001010110110011010000010;
		correct = 32'b11111011110011000000010000001011;
		#400 //1.9777045e+35 * -10.712526 = -2.1186211e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100100010011100101000001101011;
		b = 32'b01010011010110101100101011100101;
		correct = 32'b11111000001100000101001111111111;
		#400 //-1.5223296e+22 * 939706900000.0 = -1.4305436e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110011011011100000110000110110;
		b = 32'b10010101011111010111010111010000;
		correct = 32'b10001001011010111010111110011110;
		#400 //5.54248e-08 * -5.118588e-26 = -2.836967e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011100010100011001010100010000;
		b = 32'b00111110111110101101011001101100;
		correct = 32'b01011011110011010101101100011101;
		#400 //2.3596866e+17 * 0.48991716 = 1.156051e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100101000011110100100111000101;
		b = 32'b10011101101100100001111010000011;
		correct = 32'b10000011010001110110010010111110;
		#400 //1.2428267e-16 * -4.7147756e-21 = -5.859649e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000010110001110110001010110011;
		b = 32'b11011110000010100011101110100111;
		correct = 32'b00100001010101110101001101010101;
		#400 //-2.9297073e-37 * -2.4901847e+18 = 7.295512e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011110100001010111111010110001;
		b = 32'b00000111101101010110011001011010;
		correct = 32'b10100110101111010010111111100101;
		#400 //-4.80966e+18 * 2.729401e-34 = -1.3127491e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100100100101010101000001111110;
		b = 32'b01010001010011010101101110100101;
		correct = 32'b10110110011011111000110111010001;
		#400 //-6.475481e-17 * 55125365000.0 = -3.5696323e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101101100101010001000000011010;
		b = 32'b10111101000101100111110111010011;
		correct = 32'b10101011001011110100000101100110;
		#400 //1.694649e-11 * -0.03674109 = -6.226325e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101110111111110001110100111111;
		b = 32'b00011001101100001001011100111010;
		correct = 32'b11001001001011111111101011001111;
		#400 //-3.9477017e+28 * 1.8259053e-23 = -720812.94
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101101110011111111110101001111;
		b = 32'b10010101101010101101110000011100;
		correct = 32'b10000100000010101101000100001011;
		#400 //2.3645667e-11 * -6.9009725e-26 = -1.631781e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010000110001100101111100100;
		b = 32'b10100111011100110110101010101110;
		correct = 32'b00100010000100010100100100110110;
		#400 //-0.0005828722 * -3.3780856e-15 = 1.9689922e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111011011111010011011011001101;
		b = 32'b10010010001011000001110011001111;
		correct = 32'b00001110001010100011110101010000;
		#400 //-0.00386374 * -5.430914e-28 = 2.0983639e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011001010011000111001100101111;
		b = 32'b10101000100010110010111101101101;
		correct = 32'b10000010010111100101000011010101;
		#400 //1.0569814e-23 * -1.5452668e-14 = -1.6333182e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000011110101010110101010011110;
		b = 32'b01000111101101111010111110110110;
		correct = 32'b01001100000110010010000110110011;
		#400 //426.83295 * 94047.42 = 40142540.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000110011101000100000001100010;
		b = 32'b01101100100111110110110101001100;
		correct = 32'b00110011100110000001110001000101;
		#400 //4.59386e-35 * 1.5418828e+27 = 7.083194e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010011000111110101100110011;
		b = 32'b01000110110110101000110110110011;
		correct = 32'b11000001110000101001010001110001;
		#400 //-0.000869441 * 27974.85 = -24.322481
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000100101100001111000101001110;
		b = 32'b11011011001001000101000111100001;
		correct = 32'b00100000011000110010011001011100;
		#400 //-4.1599005e-36 * -4.6251923e+16 = 1.924034e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110110110011110000100011001100;
		b = 32'b00101011101010110110010110000000;
		correct = 32'b00100011000010101001110011110110;
		#400 //6.170105e-06 * 1.2178453e-12 = 7.514233e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111010110011110100101010000011;
		b = 32'b01000011001010111101001101010111;
		correct = 32'b00111110100010110010000111100110;
		#400 //0.0015815053 * 171.82555 = 0.271743
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111100111000010100010100000100;
		b = 32'b11100101100111101111110011110100;
		correct = 32'b01100011000010111110011100101111;
		#400 //-0.02749873 * -9.385001e+22 = 2.580756e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110011111110111000010111111111;
		b = 32'b10101001110110111100010110110100;
		correct = 32'b00011110010101111110110111100000;
		#400 //-1.1712472e-07 * -9.75985e-14 = 1.1431197e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110010101101000110000110110010;
		b = 32'b10111101110010111111110100000111;
		correct = 32'b00110001000011111011101111000010;
		#400 //-2.0999185e-08 * -0.099603705 = 2.0915967e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100000100101101110010001000011;
		b = 32'b11110001011000001000110001001010;
		correct = 32'b11010010100001000101101001101011;
		#400 //2.556204e-19 * -1.11190786e+30 = -284226320000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010010111101100101011010001100;
		b = 32'b00000000111110000100000001001101;
		correct = 32'b10010100011011101110000110110111;
		#400 //-529007000000.0 * 2.279827e-38 = -1.2060444e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100111100011111111001011111001;
		b = 32'b10100000100101000110000110101010;
		correct = 32'b11001000101001101101111011000101;
		#400 //1.3595609e+24 * -2.5136804e-19 = -341750.16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000011100101101001101000111111;
		b = 32'b11100100100000101110011001110011;
		correct = 32'b01101000100110100000001111001100;
		#400 //-301.20505 * -1.9317459e+22 = 5.818516e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101010110100101000110111010001;
		b = 32'b10100000100100000111011111000010;
		correct = 32'b01001011111011011010010010001010;
		#400 //-1.2727207e+26 * -2.4473798e-19 = 31148308.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011111010011101111111111110000;
		b = 32'b00010101111101000100010001101100;
		correct = 32'b10110101110001011000001101000100;
		#400 //-1.4915904e+19 * 9.8658766e-26 = -1.4715847e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101101010010001011000110011001;
		b = 32'b10001111111011011010100110010101;
		correct = 32'b00111101101110100101000101011101;
		#400 //-3.8819815e+27 * -2.3435325e-29 = 0.0909755
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110010110011100000101001000011;
		b = 32'b01100110111110101110010011010100;
		correct = 32'b11011010010010011110111000110001;
		#400 //-2.3986223e-08 * 5.9240638e+23 = -1.4209591e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001100001011011101001000100110;
		b = 32'b11100110111101111011000111110111;
		correct = 32'b01110011101010000010111010011001;
		#400 //-45566104.0 * -5.848537e+23 = 2.6649505e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011100110101010000000001101110;
		b = 32'b10110110111000010011001011111101;
		correct = 32'b11010100001110110101111111001101;
		#400 //4.7963714e+17 * -6.7114584e-06 = -3219064600000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000111010001100111110001111101;
		b = 32'b00111100001100100010010111011011;
		correct = 32'b00000100000010100001111111101001;
		#400 //1.4932448e-34 * 0.010873283 = 1.6236474e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000111101100011010010001101000;
		b = 32'b11100000101111001010011110000011;
		correct = 32'b00101001000000101110100011111010;
		#400 //-2.672863e-34 * -1.0875182e+20 = 2.9067874e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010100101111010011001011101100;
		b = 32'b01000000100010000010111111110010;
		correct = 32'b10010101110010010100110011111001;
		#400 //-1.9104208e-26 * 4.2558527 = -8.1304695e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101000001001111110001111111100;
		b = 32'b00100110000001101011001111010111;
		correct = 32'b10001110101100001010111010001111;
		#400 //-9.3197985e-15 * 4.673432e-16 = -4.3555444e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101100001011010000010000011111;
		b = 32'b10010000111011011111001110010001;
		correct = 32'b00111101101000001101000101101110;
		#400 //-8.366545e+26 * -9.385529e-29 = 0.078524455
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100101001011111011010001001000;
		b = 32'b11011010000000010001101100111110;
		correct = 32'b00111111101100010011100100010110;
		#400 //-1.5239912e-16 * -9085056000000000.0 = 1.3845546
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011111111011111000011111011011;
		b = 32'b11101110000010101011000000011001;
		correct = 32'b11001110100000011100010000000001;
		#400 //1.0144519e-19 * -1.0730455e+28 = -1088553100.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100010000111101110000110001111;
		b = 32'b10001010011101000001011100000010;
		correct = 32'b00101101000101110111110101000100;
		#400 //-7.327097e+20 * -1.17525e-32 = 8.611171e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000010101111001110110000001011;
		b = 32'b00110101110001011100111111000001;
		correct = 32'b10111001000100011111101011110110;
		#400 //-94.46102 * 1.4738108e-06 = -0.00013921768
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101001011100001000101100110101;
		b = 32'b00110110111011000001100111011011;
		correct = 32'b11100000110111011101100010100000;
		#400 //-1.8174974e+25 * 7.036358e-06 = -1.2788562e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011010001100100011001001011110;
		b = 32'b00100111001001010000100010011111;
		correct = 32'b00000001111001011100000011101110;
		#400 //3.6850224e-23 * 2.2903023e-15 = 8.4398155e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100100010010110100011110001001;
		b = 32'b11000110011011010101001000011001;
		correct = 32'b11101011001111000111001001101011;
		#400 //1.4999375e+22 * -15188.524 = -2.2781838e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001110011001001011111011101011;
		b = 32'b01111100010010001110100001110101;
		correct = 32'b01001011001100111000010011011101;
		#400 //2.8195093e-30 * 4.1726966e+36 = 11764957.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001000010000101101101001110001;
		b = 32'b11001101001010001110000101001011;
		correct = 32'b01010110000000001000101011010101;
		#400 //-199529.77 * -177083570.0 = 35333440000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100100001110110010000111001100;
		b = 32'b01010110001101110011110101111001;
		correct = 32'b10111011000001011111001000011000;
		#400 //-4.0577788e-17 * 50368663000000.0 = -0.0020438489
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011110000000110001111001100100;
		b = 32'b10101001001110110000111000111010;
		correct = 32'b10000111101111111001110011111001;
		#400 //6.941367e-21 * -4.153468e-14 = -2.8830746e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011110101111101001110100000111;
		b = 32'b11001010111101100110000110101010;
		correct = 32'b11101010001101110111001110011101;
		#400 //6.867571e+18 * -8073429.0 = -5.544485e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001111010101010100100000111110;
		b = 32'b00110110001000010111100110100111;
		correct = 32'b10000110000001101000011111001001;
		#400 //-1.0515624e-29 * 2.406168e-06 = -2.5302358e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110100100001101000001001101011;
		b = 32'b10011011011011000110001100001100;
		correct = 32'b01010000011110000110100010001011;
		#400 //-8.525549e+31 * -1.9553466e-22 = 16670404000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001100010101111010011101001100;
		b = 32'b11101110111101000110100000101001;
		correct = 32'b00111011110011011110001100110011;
		#400 //-1.6613342e-31 * -3.7820132e+28 = 0.006283188
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001011101100101010001000011100;
		b = 32'b01011110000100101110101111010110;
		correct = 32'b10101010010011010000101000001000;
		#400 //-6.880702e-32 * 2.6466977e+18 = -1.8211138e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000110000100000001011011100001;
		b = 32'b10010110011111111010000010110100;
		correct = 32'b10011101000011111110000100111110;
		#400 //9221.72 * -2.0649445e-25 = -1.904234e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101011000111110001110111010111;
		b = 32'b10101010000110100001110001011001;
		correct = 32'b00010101101111111001001100100100;
		#400 //-5.652956e-13 * -1.3687783e-13 = 7.737643e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100100100001101000011100000000;
		b = 32'b10101110110011110101100101110001;
		correct = 32'b11010011110110011110110001010011;
		#400 //1.9852732e+22 * -9.429158e-11 = -1871945500000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010110011110010110100001111010;
		b = 32'b01100010011111000110100110110100;
		correct = 32'b00111001011101011110100111010011;
		#400 //2.0147027e-25 * 1.16404905e+21 = 0.00023452127
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010000011101110001011111010000;
		b = 32'b11111100001111100101000100110100;
		correct = 32'b01001101001101111011001000001101;
		#400 //-4.8730505e-29 * -3.9527336e+36 = 192618700.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111110001001100100010111001;
		b = 32'b10010010101100101101001100100001;
		correct = 32'b00001011000010010111010111011011;
		#400 //-2.345849e-05 * -1.1285427e-27 = 2.6473905e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110001110110010110000110111101;
		b = 32'b10110001001101100100100011111111;
		correct = 32'b01100011100110101100100101111000;
		#400 //-2.152845e+30 * -2.652598e-09 = 5.710632e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011111111001011100101101110110;
		b = 32'b11011000001000001000011011100101;
		correct = 32'b00111000100100000001100001000000;
		#400 //-9.732187e-20 * -706004900000000.0 = 6.870972e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110100011001101110101111000001;
		b = 32'b11000010010001101001011111100111;
		correct = 32'b00110111001100110010001101011101;
		#400 //-2.1506186e-07 * -49.648342 = 1.0677465e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101101111101100101101011000111;
		b = 32'b01011000100000100111100101010011;
		correct = 32'b01000110111110110001110110110100;
		#400 //2.8007275e-11 * 1147660800000000.0 = 32142.852
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110001101010010111100001110;
		b = 32'b11111011111100101000010001010011;
		correct = 32'b01110010101010111010010000100010;
		#400 //-2.6998491e-06 * -2.5184394e+36 = 6.799406e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101001000111011111010001101101;
		b = 32'b10110001010010001000100001011001;
		correct = 32'b00011010111101110111011000101100;
		#400 //-3.507301e-14 * -2.9181335e-09 = 1.0234772e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100101001110111010010010110100;
		b = 32'b01100110101101101010000111000010;
		correct = 32'b01001100100001011101110110101001;
		#400 //1.6275468e-16 * 4.312273e+23 = 70184264.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110001010001100111110100001;
		b = 32'b00010001111100110000101101110111;
		correct = 32'b10001000101000000100010010100101;
		#400 //-2.5154807e-06 * 3.8345706e-28 = -9.645788e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110010111101100010110100010111;
		b = 32'b10001010110101010010001111001010;
		correct = 32'b00111110010011001111010111101111;
		#400 //-9.7520413e+30 * -2.0524616e-32 = 0.20015691
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010011000010011011001101111000;
		b = 32'b01111100011011111110010110101011;
		correct = 32'b01010000000000010000101000010111;
		#400 //1.7380316e-27 * 4.9824687e+36 = 8659688000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000010010001111010100110000001;
		b = 32'b01011111111111000101001001011100;
		correct = 32'b00100010110001001100101100010111;
		#400 //1.4668856e-37 * 3.6363392e+19 = 5.3340936e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110010001011110001000001011011;
		b = 32'b10011101111001011111111111011011;
		correct = 32'b01010000100111010100100010011000;
		#400 //-3.4674976e+30 * -6.0880344e-21 = 21110243000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011100101001011011100101111100;
		b = 32'b01001110100000111010001011101000;
		correct = 32'b11101011101010100110111011000000;
		#400 //-3.731785e+17 * 1104245800.0 = -4.120808e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000011010010001000111111100011;
		b = 32'b11111111111110101010101100111010;
		correct = 32'b11111111111110101010101100111010;
		#400 //-5.893989e-37 * nan = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001010111010011110110101011000;
		b = 32'b10111100101101100010101010110000;
		correct = 32'b01001000001001100111010110111110;
		#400 //-7665324.0 * -0.022237152 = 170454.97
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000011000100000000010000110110;
		b = 32'b11001001001110000001000111000100;
		correct = 32'b00001100110011110001101000001011;
		#400 //-4.232263e-37 * -753948.25 = 3.1909074e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000010011000111100000001001001;
		b = 32'b11101001100100110011111001101010;
		correct = 32'b10101100100000101111111011110001;
		#400 //1.6732509e-37 * -2.2250855e+25 = -3.7231264e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101001001011000001111010100010;
		b = 32'b10011011011111010101010010101100;
		correct = 32'b01000101001010100101001100110100;
		#400 //-1.3004994e+25 * -2.0955028e-22 = 2725.2002
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011101101011111000010001001011;
		b = 32'b11011001111000000001100101101110;
		correct = 32'b01111000000110011010010100110001;
		#400 //-1.5809145e+18 * -7884794400000000.0 = 1.2465186e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100101001111110001111000010011;
		b = 32'b10011000111010111001111011000110;
		correct = 32'b10111110101011111110011100100100;
		#400 //5.6407923e+22 * -6.0906396e-24 = -0.34356034
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000001111010000010111110000100;
		b = 32'b01011001100100011101001000000001;
		correct = 32'b01011100000001000100000101100010;
		#400 //29.023201 * 5130596700000000.0 = 1.4890634e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111000111100111011000101101000;
		b = 32'b01001011111111000001100000100111;
		correct = 32'b01000101011011111111100110100000;
		#400 //0.000116201874 * 33042510.0 = 3839.6016
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100000001101111011011000111100;
		b = 32'b01000111100011000011000010010011;
		correct = 32'b01101000010010010011010100001001;
		#400 //5.2951337e+19 * 71777.15 = 3.800696e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010010111011010001000000011110;
		b = 32'b10111111001011110111101100001111;
		correct = 32'b11010010101000100111111111111001;
		#400 //509088830000.0 * -0.6854715 = -348965860000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011000000000010100100010101100;
		b = 32'b11110101110101010010010000010000;
		correct = 32'b01001110010101110100011101011011;
		#400 //-1.670955e-24 * -5.403763e+32 = 902944450.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111011100000111110101000000000;
		b = 32'b00101010011100000000000001110111;
		correct = 32'b11100110011101110101011100111011;
		#400 //-1.369874e+36 * 2.1316443e-13 = -2.9200841e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111101011010111001111101000111;
		b = 32'b10101011100111110101110010010000;
		correct = 32'b01101001100100101010110100011111;
		#400 //-1.9574725e+37 * -1.1323321e-12 = 2.216509e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100111011011001010001001111111;
		b = 32'b00001001001000001111010110000011;
		correct = 32'b10110001000101001100100010000000;
		#400 //-1.117476e+24 * 1.9374738e-33 = -2.1650806e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001111100101010001000100100111;
		b = 32'b00110001101000111101000111010010;
		correct = 32'b11000001101111101100100000110010;
		#400 //-5001858600.0 * 4.767778e-09 = -23.847752
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111010010010011101001100000000;
		b = 32'b01101000000001100100000110000101;
		correct = 32'b01100010110100111011000000110011;
		#400 //0.0007698983 * 2.536023e+24 = 1.9524797e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010010011001100010000001101001;
		b = 32'b11011011011011111100100010001111;
		correct = 32'b11101110010101111000110010001100;
		#400 //247096560000.0 * -6.7493036e+16 = -1.6677297e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100100100010000110100001001011;
		b = 32'b01100110010011010100011100101111;
		correct = 32'b11001011010110101100001011100100;
		#400 //-5.915728e-17 * 2.4234956e+23 = -14336740.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010000011011011100100001010001;
		b = 32'b11100010000110000110110011110101;
		correct = 32'b11110011000011011001010000100100;
		#400 //15957313000.0 * -7.029391e+20 = -1.1217018e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110111111001001001100100000010;
		b = 32'b00111011001001100110100100001111;
		correct = 32'b00110011100101001001100100000111;
		#400 //2.7250968e-05 * 0.002539221 = 6.9196226e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110111011001101110110011111111;
		b = 32'b10001111101010000111001001010010;
		correct = 32'b01000111100101111111001010100111;
		#400 //-4.683731e+33 * -1.6610114e-29 = 77797.305
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010110010101011101010110000000;
		b = 32'b11101100110101111000011001000110;
		correct = 32'b11000011101101000000011001110111;
		#400 //1.7273372e-25 * -2.0844251e+27 = -360.0505
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111000101010100100011100101100;
		b = 32'b00001001000010101001001000111111;
		correct = 32'b01000010001110000101011101001000;
		#400 //2.7629188e+34 * 1.667991e-33 = 46.085236
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100011011010000111000101101001;
		b = 32'b00010110001110000001010011011111;
		correct = 32'b00111010001001110010010001110111;
		#400 //4.2878167e+21 * 1.4869987e-25 = 0.0006375978
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101110100110101010011100010011;
		b = 32'b00100011100111100010111101000110;
		correct = 32'b11010010101111110001111101011001;
		#400 //-2.3931336e+28 * 1.7150415e-17 = -410432340000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110101001001111100011100101011;
		b = 32'b11011110110010010100101001011010;
		correct = 32'b01010100100000111110110000011011;
		#400 //-6.2502176e-07 * -7.252252e+18 = 4532815300000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101000111111001100110010111011;
		b = 32'b00110011101001000011000010001010;
		correct = 32'b11011101001000100010001100010110;
		#400 //-9.550504e+24 * 7.645674e-08 = -7.302004e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100100101010101110100010010000;
		b = 32'b00110011100000000100001010101111;
		correct = 32'b11011000101010110100000110011010;
		#400 //-2.5221635e+22 * 5.972594e-08 = -1506386000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101000110100111101111111001111;
		b = 32'b00111100111100100001001110001101;
		correct = 32'b00100110010010000101100111000000;
		#400 //2.3522767e-14 * 0.029550338 = 6.9510573e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000010111011000011010001110000;
		b = 32'b11111111110111000101001110011100;
		correct = 32'b11111111110111000101001110011100;
		#400 //-118.10242 * nan = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011000111110001001100100011000;
		b = 32'b01110111100111001010011100010111;
		correct = 32'b11010001000110000001111110001101;
		#400 //-6.4261083e-24 * 6.354588e+33 = -40835273000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000111011100101110010101000;
		b = 32'b11101001001110010010111001100010;
		correct = 32'b01011010101011000110110000100101;
		#400 //-1.7343114e-09 * -1.3991895e+25 = 2.4266301e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010101100110001011111010010100;
		b = 32'b00101001011110011001100001000110;
		correct = 32'b10111111100101001110110000111001;
		#400 //-20993037000000.0 * 5.5421183e-14 = -1.163459
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111001111011101000110010001111;
		b = 32'b11110100011010101111001000101101;
		correct = 32'b11101110110110101110111000100110;
		#400 //0.00045499622 * -7.445736e+31 = -3.3877818e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000011000001110100101110111001;
		b = 32'b00111111011010000010000111000011;
		correct = 32'b10000010111101010101110011101111;
		#400 //-3.975986e-37 * 0.90676516 = -3.6052856e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000011100000001111011100000111;
		b = 32'b01010101001010111001000010111110;
		correct = 32'b01011001001011001101101111011001;
		#400 //257.9299 * 11789884000000.0 = 3040963800000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111000111101101100110000010100;
		b = 32'b10011101111110110101011011100110;
		correct = 32'b11010111011100100100110111011110;
		#400 //4.0045132e+34 * -6.6528998e-21 = -266416250000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101110110011111111000001110000;
		b = 32'b00110110110001110011110101010011;
		correct = 32'b10100110001000011101010110110111;
		#400 //-9.4559804e-11 * 5.9378012e-06 = -5.6147734e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111000100010100101101100000111;
		b = 32'b00000010001011100100110110101010;
		correct = 32'b00111011001111000110011110110000;
		#400 //2.2449476e+34 * 1.280579e-37 = 0.0028748326
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100110011000111010001000111110;
		b = 32'b10010100110110000000101100010101;
		correct = 32'b00111011110000000001101010111111;
		#400 //-2.687425e+23 * -2.1814797e-26 = 0.0058625634
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000010101111101110000110100101;
		b = 32'b01111000110110101001010000001000;
		correct = 32'b11111100001000101111101010000111;
		#400 //-95.44071 * 3.5466348e+34 = -3.3849336e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000110000100101011001101001;
		b = 32'b11101000110001010010000011100000;
		correct = 32'b01011010000101011010010101110100;
		#400 //-1.4139917e-09 * -7.447301e+24 = 1.0530422e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110001011010110011000001001111;
		b = 32'b01011111110101011101101111001000;
		correct = 32'b11010001110001000111100100011100;
		#400 //-3.422446e-09 * 3.082026e+19 = -105480680000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010011010110100010010110001111;
		b = 32'b11111101000001011110000010000111;
		correct = 32'b01010000111001000010100110101110;
		#400 //-2.7533986e-27 * -1.1122071e+37 = 30623494000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010101011001101111011010100011;
		b = 32'b01011001101001000010101000111011;
		correct = 32'b10101111100101000001110000011010;
		#400 //-4.6642692e-26 * 5776041000000000.0 = -2.694101e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001111101100111101101100000100;
		b = 32'b11001100010000111010101101100011;
		correct = 32'b11011100100010010111100000111101;
		#400 //6034950000.0 * -51293580.0 = -3.095542e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001101111110010001010101000000;
		b = 32'b00110100100001000111100010011110;
		correct = 32'b10000011000000001110010001010001;
		#400 //-1.5350926e-30 * 2.4674677e-07 = -3.7877914e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010000110001001110011011010110;
		b = 32'b01010001111011011000010000010101;
		correct = 32'b00100011001101101010111101001011;
		#400 //7.766403e-29 * 127515400000.0 = 9.9033595e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111000001110100001010010000111;
		b = 32'b11100001100111100001100000111101;
		correct = 32'b11011010011001011101010010010011;
		#400 //4.4364973e-05 * -3.645415e+20 = -1.6172874e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000011011110010010000010101111;
		b = 32'b11101100010011011101110100111001;
		correct = 32'b11110000010010000101011001110101;
		#400 //249.12767 * -9.9549795e+26 = -2.4800609e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100101010000100101011110011011;
		b = 32'b00010101000101100011011101001000;
		correct = 32'b00111010111001000001001010011001;
		#400 //5.7359696e+22 * 3.0335868e-26 = 0.0017400562
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010110000100110000010100101111;
		b = 32'b11010100111111000001000001111011;
		correct = 32'b01101011100100001100001010010001;
		#400 //-40412620000000.0 * -8660866000000.0 = 3.5000826e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111010001101100100101001001;
		b = 32'b00001011010001100001011101110101;
		correct = 32'b00010011000110011101000111100101;
		#400 //50889.285 * 3.815106e-32 = 1.94148e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100110111111110010100001000000;
		b = 32'b00010101101100110001110111000011;
		correct = 32'b00111101001100101000011011001111;
		#400 //6.0247297e+23 * 7.234448e-26 = 0.043585595
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001010101011010100001101000001;
		b = 32'b01101111101011011100101010000101;
		correct = 32'b11111010111010110011111100001000;
		#400 //-5677472.5 * 1.0757148e+29 = -6.107341e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010000011001100010000101100010;
		b = 32'b10111110111010100010000111100110;
		correct = 32'b01001111110100100111100011111101;
		#400 //-15443790000.0 * -0.45728987 = 7062289000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110100000011001100011100101111;
		b = 32'b00011000000110100110110001111001;
		correct = 32'b01001100101010011101011011110010;
		#400 //4.461435e+31 * 1.9958798e-24 = 89044880.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100100111100100100101011101000;
		b = 32'b00111110101101100101000001000101;
		correct = 32'b00100100001011001000110100111010;
		#400 //1.05077666e-16 * 0.35608116 = 3.7416178e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101100111000010110010111011001;
		b = 32'b00100111000111011001000110000001;
		correct = 32'b10010100100010101011101110010010;
		#400 //-6.406192e-12 * 2.1867005e-15 = -1.4008422e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001010001101001100001011100111;
		b = 32'b01011001110001010010111101000011;
		correct = 32'b11100100100010110011101101011011;
		#400 //-2961593.8 * 6937817000000000.0 = -2.0546996e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010111000001100110010001100111;
		b = 32'b00000001001010000010001101010001;
		correct = 32'b10011000101100001000100011011100;
		#400 //-147765780000000.0 * 3.0882065e-38 = -4.5633126e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110010111101111010100111110100;
		b = 32'b10011110011000010010110000111000;
		correct = 32'b01010001110110011101011100100111;
		#400 //-9.810977e+30 * -1.1920545e-20 = 116952195000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111101110111000101100111100010;
		b = 32'b01000110011011000011100100110100;
		correct = 32'b11000100110010110101010000011001;
		#400 //-0.10759331 * 15118.301 = -1626.628
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100000111010010111000101101011;
		b = 32'b11100110100001010101001110110001;
		correct = 32'b11000111111100110010100001111100;
		#400 //3.954679e-19 * -3.148093e+23 = -124496.97
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011010110001110101000101011011;
		b = 32'b01011111100000111000111010100011;
		correct = 32'b10111010110011001101101101011111;
		#400 //-8.243591e-23 * 1.8959387e+19 = -0.0015629343
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001110000011010100101110101011;
		b = 32'b01000111000010110100011110010100;
		correct = 32'b11010101100110011011111100101111;
		#400 //-592636600.0 * 35655.58 = -21130800000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110010010000000101000001100100;
		b = 32'b00110101110101010000100110000000;
		correct = 32'b11101000101000000000101000000110;
		#400 //-3.8091717e+30 * 1.5872502e-06 = -6.0461083e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101110000011100101011110000100;
		b = 32'b11111010101010011000100111101110;
		correct = 32'b11101001001111001000100011101111;
		#400 //3.236479e-11 * -4.4014786e+35 = -1.4245294e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110110011001111111000101110011;
		b = 32'b01000111110111101000010111111111;
		correct = 32'b11111110110010011001110011001001;
		#400 //-1.17609155e+33 * 113931.99 = -1.3399445e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010111101111010111110010011111;
		b = 32'b01110111000001100111110001011110;
		correct = 32'b11001111010001110001011010010010;
		#400 //-1.2245298e-24 * 2.7276963e+33 = -3340145200.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101101100111011111001011101101;
		b = 32'b00100101101100001111001101001010;
		correct = 32'b00010011110110100101101000111100;
		#400 //1.7956714e-11 * 3.0695992e-16 = 5.5119915e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100001001101111101011101000011;
		b = 32'b01111110011001010111101001110011;
		correct = 32'b01100000001001001100101101111110;
		#400 //6.228771e-19 * 7.625725e+37 = 4.7498894e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000011011011001000101001001001;
		b = 32'b10011011100101011111100001111101;
		correct = 32'b10011111100010101001001000010110;
		#400 //236.54018 * -2.4810564e-22 = -5.868695e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000000110010000000010000100001;
		b = 32'b11101001100111111100000100110010;
		correct = 32'b00101010111110011010001100000101;
		#400 //-1.836858e-38 * -2.4141443e+25 = 4.4344403e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000010111000111010101110101111;
		b = 32'b00011011110011100001010011110110;
		correct = 32'b00011111001101110100011011001011;
		#400 //113.83532 * 3.4093387e-22 = 3.8810316e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111001001111011110001000110110;
		b = 32'b00000101101010111010011101101101;
		correct = 32'b00111111011111101010010010010011;
		#400 //6.1620763e+34 * 1.6142265e-35 = 0.9946987
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000110001011100011000111000011;
		b = 32'b11110011010101110011011001011011;
		correct = 32'b11111010000100100111000011000111;
		#400 //11148.44 * -1.7050877e+31 = -1.9009068e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000011110100000111000111111001;
		b = 32'b10000000000000100100111010110011;
		correct = 32'b00000001111100000111110000110110;
		#400 //-416.8904 * -2.11903e-40 = 8.834031e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101001111111000110011010001011;
		b = 32'b11010100101010101010011001100100;
		correct = 32'b10111111001010000100000000100101;
		#400 //1.12088365e-13 * -5863488000000.0 = -0.65722877
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010000001110110010111000101100;
		b = 32'b01001001000100101011001110100100;
		correct = 32'b10011001110101101000011101011101;
		#400 //-3.6914817e-29 * 600890.25 = -2.2181754e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110100011100011011000001111101;
		b = 32'b10000010010011100100101001001110;
		correct = 32'b10110111010000101100001000101011;
		#400 //7.659443e+31 * -1.5155814e-37 = -1.1608509e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101010111000110001000000100001;
		b = 32'b11101010001000011110011010110111;
		correct = 32'b11010101100011111001100111001000;
		#400 //4.0334492e-13 * -4.8931644e+25 = -19736330000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111101000011101010111101101000;
		b = 32'b10101001101011111100110001101001;
		correct = 32'b11100111010000111111011110101101;
		#400 //1.1853821e+37 * -7.807021e-14 = -9.254303e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110001101111101001111011000001;
		b = 32'b10111011100101101110101000001111;
		correct = 32'b11101101111000001011111010011011;
		#400 //1.8878104e+30 * -0.0046055387 = -8.694384e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000101110010111111001011010010;
		b = 32'b00000010101001101111100000101110;
		correct = 32'b10001001000001010000010100101100;
		#400 //-6526.3525 * 2.4533956e-37 = -1.6011724e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000010000001101000100100110011;
		b = 32'b01111101101010010111011001111011;
		correct = 32'b11000000001100100001110110101101;
		#400 //-9.884139e-38 * 2.815684e+37 = -2.7830613
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000000010001010010011101111000;
		b = 32'b10110110110011101011011001100111;
		correct = 32'b00110111100111110011001000111100;
		#400 //-3.080534 * -6.160513e-06 = 1.897767e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111110101100101001011001110000;
		b = 32'b10011111000011011010001110111111;
		correct = 32'b00011110010001011001111000101101;
		#400 //-0.348804 * -2.999336e-20 = 1.0461803e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101001010111001011111010000100;
		b = 32'b11111111110110100100001101011110;
		correct = 32'b11111111110110100100001101011110;
		#400 //4.901506e-14 * nan = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011000110110111000111111011000;
		b = 32'b11011100001000011011001001000110;
		correct = 32'b00110101100010101010111001011101;
		#400 //-5.675542e-24 * -1.8205394e+17 = 1.0332548e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010110011110001000111000011001;
		b = 32'b01001010111100001100011000010011;
		correct = 32'b10100001111010011100010110001000;
		#400 //-2.0078119e-25 * 7889673.5 = -1.584098e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110100101001101101101110101010;
		b = 32'b11010100100111101110111010101010;
		correct = 32'b11001001110011110010111001000100;
		#400 //3.1079736e-07 * -5460871600000.0 = -1697224.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010011000010010111111100011111;
		b = 32'b11011100110010000001111100100010;
		correct = 32'b10110000010101101111100000010010;
		#400 //1.7354507e-27 * -4.506338e+17 = -7.8205276e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101010000011010000001110011011;
		b = 32'b11011100110110101101011101001101;
		correct = 32'b01000111011100010001011101010101;
		#400 //-1.2524567e-13 * -4.9278617e+17 = 61719.332
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100110001000101000101001010111;
		b = 32'b11000101101101111011000110000110;
		correct = 32'b00101100011010010100001100110110;
		#400 //-5.6392526e-16 * -5878.1904 = 3.31486e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001100011010001001101100110100;
		b = 32'b11101010111111001001001000001100;
		correct = 32'b11110111111001010111110101111011;
		#400 //60976336.0 * -1.526695e+26 = -9.309227e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010001000100000000010100110111;
		b = 32'b01110010111100011101010101110100;
		correct = 32'b01000100100010000000110011111110;
		#400 //1.1361204e-28 * 9.580024e+30 = 1088.406
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101101000010101110101110101010;
		b = 32'b11001111100001100111101011100100;
		correct = 32'b10111101000100011111010000010110;
		#400 //7.89672e-12 * -4512401400.0 = -0.03563317
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000111110110000101011101011101;
		b = 32'b00011110000010110010110100110110;
		correct = 32'b10100110011010110011101101001001;
		#400 //-110766.73 * 7.367948e-21 = -8.161235e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110110000100000101010100011011;
		b = 32'b10001111000110101011001110001010;
		correct = 32'b01000101101011100111000011010111;
		#400 //-7.318524e+32 * -7.627364e-30 = 5582.105
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010001000001111110110110011110;
		b = 32'b01111011111100010111000001110100;
		correct = 32'b11001101100000000011001001100111;
		#400 //-1.0722844e-28 * 2.5072487e+36 = -268848350.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111111010110100010011011000;
		b = 32'b11100111010101111010110101000001;
		correct = 32'b01011111110001100011011000001011;
		#400 //-2.8046241e-05 * -1.0185048e+24 = 2.856523e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011010001001000010111011011101;
		b = 32'b01011111111111010110010100010111;
		correct = 32'b11111010101000101000001100100110;
		#400 //-1.1553356e+16 * 3.6518051e+19 = -4.2190605e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011111111110010101011110011001;
		b = 32'b00110011110110001010010101000010;
		correct = 32'b01010100010100110000001011011111;
		#400 //3.5933995e+19 * 1.0088344e-07 = 3625145000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000100010110010110011110001011;
		b = 32'b11001111101011001011111100000100;
		correct = 32'b10010100100100101011001111001001;
		#400 //2.5555772e-36 * -5796399000.0 = -1.4813145e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011111010100000011100001011010;
		b = 32'b10000110010011000111010111110010;
		correct = 32'b10100110001001100100110011010110;
		#400 //1.5003841e+19 * -3.8454788e-35 = -5.769695e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111000111010000000111101001101;
		b = 32'b01011010011011100111001100000000;
		correct = 32'b11010011110110000010011001111000;
		#400 //-0.00011065472 * 1.6779372e+16 = -1856716700000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101010101011001001101100000110;
		b = 32'b11001011011111100000100001110011;
		correct = 32'b01110110101010110100011110000010;
		#400 //-1.0433366e+26 * -16648307.0 = 1.7369787e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111110111110101011100110111010;
		b = 32'b10010001111001010100010010100100;
		correct = 32'b11010001011000001000101101011101;
		#400 //1.6663567e+38 * -3.6172133e-28 = -60275675000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100001100011100110110101111;
		b = 32'b00010001000010000101000111011100;
		correct = 32'b00010101101111010101110001000000;
		#400 //711.2138 * 1.0753733e-28 = 7.6482037e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000100001000000111111001010111;
		b = 32'b11111000110101010110100111110010;
		correct = 32'b01111101100001011100101110001010;
		#400 //-641.97406 * -3.4628377e+34 = 2.223052e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011100011111001110001110111001;
		b = 32'b00010101001111110100011110011100;
		correct = 32'b00110010001111001111010010100100;
		#400 //2.8472831e+17 * 3.8628633e-26 = 1.0998665e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101011010011011110110101001001;
		b = 32'b10010010111000110011101100010110;
		correct = 32'b10111110101101101100100011101111;
		#400 //2.4895034e+26 * -1.434028e-27 = -0.35700175
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111110011101110101000010110111;
		b = 32'b00001000000101000111111010000110;
		correct = 32'b11000111000011110111010011100101;
		#400 //-8.2184603e+37 * 4.4685858e-34 = -36724.895
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010001101001010010111111111000;
		b = 32'b10000011000001110000000101000101;
		correct = 32'b00010101001011100011101000111011;
		#400 //-88684300000.0 * -3.967439e-37 = 3.5184956e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000001100100000011101111111000;
		b = 32'b01101110010011000001001101101000;
		correct = 32'b00110000011001011111010101110001;
		#400 //5.2983297e-38 * 1.5789601e+28 = 8.365851e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110001010111011011101100100001;
		b = 32'b01101110100001010010011110110111;
		correct = 32'b11100000011001101010100100111100;
		#400 //-3.2266103e-09 * 2.060476e+28 = -6.6483527e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110101101001101011100111001110;
		b = 32'b10101010001110000101101010001001;
		correct = 32'b10100000011100000010000100000101;
		#400 //1.242204e-06 * -1.6373894e-13 = -2.0339716e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000010011000000000010011001000;
		b = 32'b11001111100001111111001100001000;
		correct = 32'b11010010011011011110111001100010;
		#400 //56.00467 * -4561703000.0 = -255476660000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010101011110101001011010101100;
		b = 32'b10000010001110000100000001111101;
		correct = 32'b00011000001101000101101101101100;
		#400 //-17220315000000.0 * -1.3536692e-37 = 2.331061e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010001000010110100001011011011;
		b = 32'b00110111010001101000001000111001;
		correct = 32'b00001000110101111111100100011001;
		#400 //1.0985768e-28 * 1.18320395e-05 = 1.2998404e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010000000011011010100101011100;
		b = 32'b00010011110100011101101010101101;
		correct = 32'b00100100011010000100000010001100;
		#400 //9506746000.0 * 5.297465e-27 = 5.0361654e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111100110100100010010110111111;
		b = 32'b00001101110000111101010010010010;
		correct = 32'b01001011001000001100000101000000;
		#400 //8.7291834e+36 * 1.2068977e-30 = 10535232.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111110101110011100000110010110;
		b = 32'b00100011010100100011100001111101;
		correct = 32'b11100010100110001000100111001010;
		#400 //-1.2345617e+38 * 1.1396085e-17 = -1.4069169e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101010100010110000000110000011;
		b = 32'b00110110000100101000001111100010;
		correct = 32'b10100001000111110001110011110010;
		#400 //-2.469241e-13 * 2.1832461e-06 = -5.3909604e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110100000000011100001011010000;
		b = 32'b01000110000100111101011111000011;
		correct = 32'b01111010100101011110000001110110;
		#400 //4.11229e+31 * 9461.94 = 3.8910242e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111110000000011110011001111011;
		b = 32'b10111110010000111011100100001001;
		correct = 32'b00111100110001101010000011101000;
		#400 //-0.12685578 * -0.19113554 = 0.024246648
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101111010111110010000000100001;
		b = 32'b10101111101010001110100010101011;
		correct = 32'b11011111100100110011011111100000;
		#400 //6.9054e+28 * -3.0724343e-10 = -2.1216387e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001110000000000000111010101101;
		b = 32'b00011000101011111111000111101011;
		correct = 32'b00100111001100000000011000010111;
		#400 //537111360.0 * 4.5480714e-24 = 2.4428208e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101110000000110010000100101101;
		b = 32'b10010100101000100100011101111111;
		correct = 32'b11000011001001100011111100111011;
		#400 //1.0145661e+28 * -1.638602e-26 = -166.247
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010111100110110101010010101011;
		b = 32'b11010001100110111001010111010100;
		correct = 32'b10101001101111001100111001011001;
		#400 //1.0038013e-24 * -83529200000.0 = -8.384673e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010100011011001011111001110101;
		b = 32'b10001001111011111101110000100011;
		correct = 32'b00011110110111011101000101100011;
		#400 //-4067230500000.0 * -5.7744173e-33 = 2.3485885e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000110011011111111101001101110;
		b = 32'b01101110110000110101010100010101;
		correct = 32'b00110101101101110001101110000100;
		#400 //4.513489e-35 * 3.0226217e+28 = 1.3642571e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111001100000101000001110000101;
		b = 32'b11101010101001011110001011110100;
		correct = 32'b11100100101010010010010011110010;
		#400 //0.00024893522 * -1.0027226e+26 = -2.4961296e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000110101010011010000010010001;
		b = 32'b01101110010101101110111010010011;
		correct = 32'b11110101100011100110101001001110;
		#400 //-21712.283 * 1.6629553e+28 = -3.6106556e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000001001111000110001110001011;
		b = 32'b01011111110000001010011101100010;
		correct = 32'b11100001100011011100010111010101;
		#400 //-11.7743025 * 2.7764344e+19 = -3.2690578e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001011010001111000011000100001;
		b = 32'b11110111111111101101011111110000;
		correct = 32'b01000011110001101001111101100001;
		#400 //-3.8426913e-32 * -1.0337681e+34 = 397.24515
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010001011110000011011010111111;
		b = 32'b11110101010001101101111100111110;
		correct = 32'b11000111010000001101001011001100;
		#400 //1.958062e-28 * -2.5210026e+32 = -49362.797
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100010111010101000100100010010;
		b = 32'b11111111000100011001000010111101;
		correct = 32'b01100010100001010101110000111101;
		#400 //-6.3570956e-18 * -1.9348958e+38 = 1.2300317e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001101010101011001010101011101;
		b = 32'b10011011111000111101001100001101;
		correct = 32'b00101001101111100001001110000110;
		#400 //-223958480.0 * -3.7690388e-22 = 8.441082e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011010100101101011011101101011;
		b = 32'b11101010101011111011101001111001;
		correct = 32'b11000101110011101110101001010101;
		#400 //6.2334874e-23 * -1.06221305e+26 = -6621.2915
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110100000111000110000100110100;
		b = 32'b01111111010111111000000100110001;
		correct = 32'b01110100000010001000011110010111;
		#400 //1.4563994e-07 * 2.9708864e+38 = 4.3267973e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010111000000101110110001101110;
		b = 32'b11001001111010110110010100100000;
		correct = 32'b10100001011100001100010110000001;
		#400 //4.230368e-25 * -1928356.0 = -8.1576557e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101110100100010001010001000110;
		b = 32'b11110000110011011110000001001100;
		correct = 32'b01011111111010010101100010110010;
		#400 //-6.597438e-11 * -5.097247e+29 = 3.362877e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110000101101110010001010110110;
		b = 32'b00110010000110010001011110000111;
		correct = 32'b11100011010110110000100100100111;
		#400 //-4.5342176e+29 * 8.911122e-09 = -4.0404964e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110110110110010110111001110101;
		b = 32'b11000000000011100011010111001001;
		correct = 32'b10110111011100011001000111100111;
		#400 //6.479963e-06 * -2.2220328 = -1.439869e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111010111110011110111100000000;
		b = 32'b00011001100111101010000101100110;
		correct = 32'b11010101000110101101111100010101;
		#400 //-6.488647e+35 * 1.6402005e-23 = -10642683000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111000011100101010111001110;
		b = 32'b10011001001010001100101000110000;
		correct = 32'b00010000101110111011000101110011;
		#400 //-8.4838375e-06 * -8.726228e-24 = 7.40319e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100110110100110011100111000011;
		b = 32'b01011101100011101011100001000111;
		correct = 32'b11000100111010111000010000101101;
		#400 //-1.4656722e-15 * 1.285506e+18 = -1884.1305
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111011101100001100110000101000;
		b = 32'b10100011001110111100111000010000;
		correct = 32'b11011111100000011011001101110001;
		#400 //1.83597e+36 * -1.0180926e-17 = -1.8691876e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110101100100011101101001101000;
		b = 32'b10010000110110010001001100110111;
		correct = 32'b10000110111101110101101000101001;
		#400 //1.0866906e-06 * -8.5621013e-29 = -9.304355e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001000111000100101001010101110;
		b = 32'b10010101100010000110101001101001;
		correct = 32'b10011110111100010011001111111111;
		#400 //463509.44 * -5.509785e-26 = -2.5538373e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011111001000000110010000110010;
		b = 32'b11111000010011010011101001011011;
		correct = 32'b11011000000000001001010011001100;
		#400 //3.3964198e-20 * -1.665007e+34 = -565506260000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000010011111100010010101000001;
		b = 32'b11011000000001100101010111001100;
		correct = 32'b00011011000001010101110010101101;
		#400 //-1.8671664e-37 * -590812200000000.0 = 1.1031447e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001001010100010101111001010101;
		b = 32'b10100111001111010011001110011000;
		correct = 32'b00110001000110101011110011010111;
		#400 //-857573.3 * -2.6256988e-15 = 2.2517292e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100110101011111001101100110100;
		b = 32'b00011011111110000110011111100000;
		correct = 32'b11000011001010100110010110011011;
		#400 //-4.1463856e+23 * 4.1095286e-22 = -170.3969
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100010000111100010111010010100;
		b = 32'b00101110011101010000010001001111;
		correct = 32'b11010001000101110110010100111101;
		#400 //-7.294855e+20 * 5.5710377e-11 = -40639910000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110000000011010000110100011100;
		b = 32'b10010110111101111100000100011100;
		correct = 32'b11000111100010001000001000001100;
		#400 //1.7461294e+29 * -4.0026871e-25 = -69892.09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101101000010100110110100111110;
		b = 32'b11001111100110101100010110000000;
		correct = 32'b11111101001001110110000100000101;
		#400 //2.6775623e+27 * -5193269000.0 = -1.3905302e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101100000000010011110110011100;
		b = 32'b10001011110011101001111011000110;
		correct = 32'b00111000010100001001111101110111;
		#400 //-6.249695e+26 * -7.958721e-32 = 4.9739578e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010000011010101010010110001110;
		b = 32'b01011000100111010000100100000001;
		correct = 32'b00101001100011111110111111001001;
		#400 //4.6275902e-29 * 1381296000000000.0 = 6.392072e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110101101010010010011100010101;
		b = 32'b00110101000000110100110111010111;
		correct = 32'b01101011001011011000010011011101;
		#400 //4.2885295e+32 * 4.8914575e-07 = 2.097716e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111011101100001001011110111011;
		b = 32'b00001001100110011001010111100010;
		correct = 32'b00000101110100111110010000100110;
		#400 //0.0053891814 * 3.697436e-33 = 1.9926153e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111010011011111001011001000001;
		b = 32'b00010011011110000101110100100010;
		correct = 32'b01001110011010000111000010111000;
		#400 //3.1100162e+35 * 3.1347919e-27 = 974925300.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101001100011010000110010000101;
		b = 32'b10110101101001111010111010110110;
		correct = 32'b01011111101110001100011011011011;
		#400 //-2.1314708e+25 * -1.2493317e-06 = 2.662914e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011101110110111010101001001000;
		b = 32'b00110101110100000001011010011000;
		correct = 32'b00010100001100101000110110111110;
		#400 //5.8144884e-21 * 1.5503783e-06 = 9.014657e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111111111000101100011000011110;
		b = 32'b01110100100111010111011001110010;
		correct = 32'b11110101000010110111110001101101;
		#400 //-1.771671 * 9.980383e+31 = -1.7681956e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100000101101101010010000111000;
		b = 32'b11101110111100000010110111000001;
		correct = 32'b11010000001010110101101010011001;
		#400 //3.094067e-19 * -3.7165858e+28 = -11499365000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111001111000111010101000100000;
		b = 32'b10111011010111100111000011011101;
		correct = 32'b10110101110001011101000111100111;
		#400 //0.00043423567 * -0.0033941783 = -1.4738733e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100111000111000001101000100001;
		b = 32'b11000101001001011111100001100011;
		correct = 32'b11101100110010100110100010011010;
		#400 //7.371712e+23 * -2655.5242 = -1.9575759e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000010110010101011011001110101;
		b = 32'b11110010010101001110000000010110;
		correct = 32'b10110101101010001001000010001010;
		#400 //2.9785958e-37 * -4.2164304e+30 = -1.2559042e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001101111101100010100110011101;
		b = 32'b01010110010010001110110100001101;
		correct = 32'b01100100110000010011010001110100;
		#400 //516240300.0 * 55230113000000.0 = 2.851201e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111001011101101111110101111010;
		b = 32'b00110100101000101111001100100100;
		correct = 32'b10101110100111010011011011111101;
		#400 //-0.00023554816 * 3.035176e-07 = -7.149301e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001011100011101110111101101000;
		b = 32'b11011110100110101001100100111010;
		correct = 32'b10101010101011001010001100100100;
		#400 //5.505663e-32 * -5.5699995e+18 = -3.066654e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110100111010101011101010011;
		b = 32'b01100000011101111100100010011100;
		correct = 32'b01011111100110000100101010001101;
		#400 //0.30730686 * 7.141877e+19 = 2.1947477e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011000000010011001000001000111;
		b = 32'b01001001110111111011101000100001;
		correct = 32'b10100010011100000111000101100101;
		#400 //-1.7779676e-24 * 1832772.1 = -3.2586096e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110101000101110110110110101011;
		b = 32'b10100010000000111000101000101110;
		correct = 32'b00010111100110111001110110110110;
		#400 //-5.641147e-07 * -1.7826962e-18 = 1.0056452e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000001101101101101101101000101;
		b = 32'b01111111000001100100001011111110;
		correct = 32'b11000001001111111100110101000000;
		#400 //-6.717088e-38 * 1.784644e+38 = -11.98761
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011100101010001011111111101100;
		b = 32'b10101100100101010111000001100100;
		correct = 32'b00001001110001010000001110010100;
		#400 //-1.1166918e-21 * -4.2473126e-12 = 4.742939e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011111000101010111100100101000;
		b = 32'b00101001010011010100010000110000;
		correct = 32'b01001000111011111011001110101010;
		#400 //1.0770684e+19 * 4.5578287e-14 = 490909.3
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001001111000110110110101110000;
		b = 32'b11111101001100000011110011001001;
		correct = 32'b01000111100111001001000100111101;
		#400 //-5.4751177e-33 * -1.4641234e+37 = 80162.48
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001011011100001001111010110110;
		b = 32'b11011011010110110100100011010011;
		correct = 32'b00100111010011100001110000111001;
		#400 //-4.634172e-32 * -6.172309e+16 = 2.8603542e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110100110011001001011111111111;
		b = 32'b00011010111110110110011010011001;
		correct = 32'b11010000010010001110101100000110;
		#400 //-1.2967669e+32 * 1.0397692e-22 = -13483383000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101101010100100111101010100110;
		b = 32'b00111000110101001011011000001100;
		correct = 32'b00100110101011101110001100111111;
		#400 //1.1964351e-11 * 0.000101428566 = 1.2135271e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111111101001101001100110011111;
		b = 32'b11111001011110110011011010101001;
		correct = 32'b11111001101000110111110000110001;
		#400 //1.3015631 * -8.1523447e+34 = -1.0610791e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001100000101110001011100000000;
		b = 32'b00111010111000001110001100001101;
		correct = 32'b10000111100001001011101000100001;
		#400 //-1.1639538e-31 * 0.001715751 = -1.997055e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111011011101011000011110111100;
		b = 32'b10110101111000011111101000011011;
		correct = 32'b00110001110110001011110000101101;
		#400 //-0.0037464937 * -1.6836597e-06 = 6.3078205e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101001000010110101001011111111;
		b = 32'b10101010100001001010010110000111;
		correct = 32'b11010100000100000110000111000011;
		#400 //1.0527039e+25 * -2.3562768e-13 = -2480461800000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010100010001001010100001110110;
		b = 32'b00010011101111100111001110001101;
		correct = 32'b00101000100100100100110111001100;
		#400 //3378559600000.0 * 4.8076685e-27 = 1.6242995e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111011111100101110100110110101;
		b = 32'b00101110010100001010010100010101;
		correct = 32'b10101010110001011111101010001000;
		#400 //-0.007413114 * 4.7440347e-11 = -3.516807e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100011000111010000011111010;
		b = 32'b10001111100001000110111010001011;
		correct = 32'b10010100011010111000001010010111;
		#400 //910.51526 * -1.3058785e-29 = -1.1890222e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111001111110001100010000111111;
		b = 32'b00101011000110100100110110110100;
		correct = 32'b11100101100101011111000110010000;
		#400 //-1.6145875e+35 * 5.4819625e-13 = -8.851108e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100011100011111100101000011100;
		b = 32'b00000111111010000011010101011110;
		correct = 32'b10101100000000100110110100100011;
		#400 //-5.304896e+21 * 3.4938847e-34 = -1.8534694e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110101011001100000101011001001;
		b = 32'b10011100000111010001001100101100;
		correct = 32'b10010010000011010010010111011000;
		#400 //8.569737e-07 * -5.197172e-22 = -4.45384e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101100100000110110010010111011;
		b = 32'b10101001101010100011011110100001;
		correct = 32'b01010110101011101011101011100011;
		#400 //-1.2707597e+27 * -7.5591666e-14 = 96058850000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101110111111110011010101100110;
		b = 32'b10101100001010000101110100111010;
		correct = 32'b11011011101001111101011111111011;
		#400 //3.9491616e+28 * -2.3925987e-12 = -9.448759e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101110011100010110100011111000;
		b = 32'b01011100100101010000000000110110;
		correct = 32'b01001011100011001000001001001011;
		#400 //5.4890287e-11 * 3.3552003e+17 = 18416790.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111101100111001100011011101110;
		b = 32'b11001100100010111000101010101011;
		correct = 32'b11001010101010101110100111011110;
		#400 //0.0765513 * -73160024.0 = -5600495.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000101001101000000100101001001;
		b = 32'b00100001010110111010100101100101;
		correct = 32'b10100111000110100111101100010011;
		#400 //-2880.5803 * 7.442428e-19 = -2.1438512e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011101001001110000110100010011;
		b = 32'b01101010110000001100101010111011;
		correct = 32'b01001000011110111001110000110001;
		#400 //2.2109025e-21 * 1.1653556e+26 = 257648.77
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110101000011011001110000111111;
		b = 32'b00011101100011110010001100110111;
		correct = 32'b00010011000111100101101110000100;
		#400 //5.275396e-07 * 3.7888196e-21 = 1.9987524e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101001000001101001100010001010;
		b = 32'b00011100101011111000001111110001;
		correct = 32'b00000110001110001000111101001010;
		#400 //2.9886284e-14 * 1.1614635e-21 = 3.4711826e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111010111100110001001010010011;
		b = 32'b00000010110101111001001010111010;
		correct = 32'b00111110010011001010111111101011;
		#400 //6.3105243e+35 * 3.1675628e-37 = 0.19988982
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110011001100111000101010100111;
		b = 32'b10110010100011100100011001110111;
		correct = 32'b10100110010001111001000010101000;
		#400 //4.180279e-08 * -1.656302e-08 = -6.923804e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011110001101011001000111000111;
		b = 32'b01000011100001110110000010001010;
		correct = 32'b10100010010000000000100010110001;
		#400 //-9.612206e-21 * 270.7542 = -2.6025453e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111101110101000100001101100111;
		b = 32'b10010010011110011111000010000001;
		correct = 32'b00010000110011110011110011111001;
		#400 //-0.103644185 * -7.886699e-28 = 8.1741047e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010010000010110100001001001111;
		b = 32'b10000000111111101100010001010100;
		correct = 32'b00010011100010101001011010010111;
		#400 //-149528230000.0 * -2.3396645e-38 = 3.498459e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101111101110111111000001111111;
		b = 32'b00011101101001100101101111001111;
		correct = 32'b01001101111101000100001010110010;
		#400 //1.1632888e+29 * 4.403476e-21 = 512251460.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101001001001110111000011101001;
		b = 32'b10000000000000110001111000001111;
		correct = 32'b00100111100000100111111011110001;
		#400 //-1.2651488e+25 * -2.8629e-40 = 3.621988e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000101101001100001101001111100;
		b = 32'b11001111010001011101100100010001;
		correct = 32'b01010101100000000101111100111001;
		#400 //-5315.3105 * -3319337200.0 = 17643308000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111010011011111100001111011101;
		b = 32'b00110010100101110001100100100100;
		correct = 32'b00101101100011011000010000010011;
		#400 //0.00091463124 * 1.7590146e-08 = 1.6088497e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101101101110110010100000001111;
		b = 32'b11111000101110000111101111111011;
		correct = 32'b11100111000001101101111101101111;
		#400 //2.1277228e-11 * -2.993429e+34 = -6.369187e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000010111011010001001010110000;
		b = 32'b10110100101000011011100110000100;
		correct = 32'b00111000000101011100010010001101;
		#400 //-118.5365 * -3.0123567e-07 = 3.570742e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001110101101100101001010110001;
		b = 32'b01101111011101011110011000010011;
		correct = 32'b00111110101011110010000011111111;
		#400 //4.4946093e-30 * 7.610197e+28 = 0.34204862
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110000100001000110101000101000;
		b = 32'b00110110000111011100000011101110;
		correct = 32'b00100111001000110011000111001011;
		#400 //9.634435e-10 * 2.3507123e-06 = 2.2647787e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010111000101011011101110100111;
		b = 32'b00110000011110111100001100101101;
		correct = 32'b11001000000100110100000100100101;
		#400 //-164633200000000.0 * 9.159063e-10 = -150788.58
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010000011000001001000100111001;
		b = 32'b11001000000111010100100001110011;
		correct = 32'b00011001000010011111100010011110;
		#400 //-4.4288086e-29 * -161057.8 = 7.132942e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011111111100010011110111001110;
		b = 32'b01000000111000011010111100000001;
		correct = 32'b10100001010101001010110000111100;
		#400 //-1.0216972e-19 * 7.052613 = -7.2056344e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110001110010101000110011000001;
		b = 32'b10111110010000100011001000110111;
		correct = 32'b11110000100110011010011001100101;
		#400 //2.0059563e+30 * -0.18964468 = -3.8041892e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101000111010101111110100110000;
		b = 32'b00010101001111001001101101011100;
		correct = 32'b10111110101011010010000010001011;
		#400 //-8.877634e+24 * 3.8088855e-26 = -0.3381389
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000011010110111001111100100011;
		b = 32'b11000110100111000111101000101000;
		correct = 32'b10001010100001100011110111000101;
		#400 //6.4540996e-37 * -20029.078 = -1.2926966e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111101111011101110101010110101;
		b = 32'b10011000101111110001010110111110;
		correct = 32'b11010111001100100101010101101000;
		#400 //3.9696866e+37 * -4.9394297e-24 = -196079890000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100010111101110100010101010000;
		b = 32'b01000001000010001101011010100110;
		correct = 32'b00100100100001000010110000100111;
		#400 //6.702287e-18 * 8.552404 = 5.732067e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101011110100001100010011101010;
		b = 32'b00110101000110100001000000101101;
		correct = 32'b10100001011110110100011101001100;
		#400 //-1.4833944e-12 * 5.739301e-07 = -8.513647e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001011100100000001111010010001;
		b = 32'b10111000110100011011111010111101;
		correct = 32'b11000100111011000010100010101011;
		#400 //18890018.0 * -0.000100014244 = -1889.2709
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111011111110000000100100100011;
		b = 32'b01011000011011111000010001100111;
		correct = 32'b11010100111010000001000011010000;
		#400 //-0.0075694486 * 1053407800000000.0 = -7973716000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110111000111011010111110111100;
		b = 32'b10110101111111010110011100000001;
		correct = 32'b11101101100111000001011000011111;
		#400 //3.1982614e+33 * -1.8879947e-06 = -6.0383005e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001111110101000010011100101011;
		b = 32'b11010101001001100111100000011011;
		correct = 32'b10100101100010011111010011101111;
		#400 //2.0919901e-29 * -11439674000000.0 = -2.3931685e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001110010111110011111011110110;
		b = 32'b11110011101101001101111101110111;
		correct = 32'b01000010100111011011101100100101;
		#400 //-2.7517187e-30 * -2.8660457e+31 = 78.86552
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000010101110001110100011100110;
		b = 32'b01101010101100111010011000110111;
		correct = 32'b00101110000000011100001011101000;
		#400 //2.7170047e-37 * 1.0859132e+26 = 2.9504316e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010000111110000001000000101110;
		b = 32'b00000101011100000110010101101001;
		correct = 32'b00010110111010001111000101101111;
		#400 //33294480000.0 * 1.1303372e-35 = 3.7633988e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100011000010000100100000010000;
		b = 32'b10011111000001111100111010101000;
		correct = 32'b00000010100100001001100000001000;
		#400 //-7.387835e-18 * -2.8758304e-20 = 2.124616e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100110011010011100011110001000;
		b = 32'b11010011010111101101010010100010;
		correct = 32'b01111010010010110111110100110101;
		#400 //-2.7599802e+23 * -957050100000.0 = 2.6414394e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011111001010011000111101101001;
		b = 32'b11100111000001000011000010000001;
		correct = 32'b01000110101011110001110000100101;
		#400 //-3.5905768e-20 * -6.242471e+23 = 22414.072
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111011011001010101011100111101;
		b = 32'b01010001110110011111011001101111;
		correct = 32'b01001101110000110100001110111000;
		#400 //0.0034994625 * 117017800000.0 = 409499400.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101001010101101000011100111000;
		b = 32'b01110100100011110001001010111110;
		correct = 32'b11011110011011111100101001111010;
		#400 //-4.763483e-14 * 9.068342e+31 = -4.3196893e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101011111101010111101100111111;
		b = 32'b00111101101101001010110011001001;
		correct = 32'b10101010001011010100000001011000;
		#400 //-1.7442505e-12 * 0.08822019 = -1.538781e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001010100000011000111011001010;
		b = 32'b10100110011011010100111101110101;
		correct = 32'b00110001011100000011001011001111;
		#400 //-4245349.0 * -8.2333577e-16 = 3.4953478e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111110100010001000101010000011;
		b = 32'b11001010111110111101110011111001;
		correct = 32'b01001010000001100101010110101010;
		#400 //-0.26668176 * -8253052.5 = 2200938.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100000110110110111101101101001;
		b = 32'b00100011001110101111001110110101;
		correct = 32'b10000100101000000100100010011100;
		#400 //-3.718171e-19 * 1.0134687e-17 = -3.76825e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001011110110011011001010001011;
		b = 32'b01100010011100001111011101101001;
		correct = 32'b01101110110011001110100111000111;
		#400 //28534038.0 * 1.1112616e+21 = 3.170878e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100001110110001000010100001011;
		b = 32'b01011000101101111010011100010110;
		correct = 32'b00111011000110110101010001101100;
		#400 //1.4671946e-18 * 1615426000000000.0 = 0.0023701442
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010100011110111100100001011110;
		b = 32'b10100001111010010100000000011011;
		correct = 32'b00110110111001010110100001101010;
		#400 //-4325593600000.0 * -1.5805663e-18 = 6.836887e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100001011001010000001010111001;
		b = 32'b00010000110110001110000101110011;
		correct = 32'b00110010110000100000001111111010;
		#400 //2.6403129e+20 * 8.554434e-29 = 2.258638e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001010100100000100011110010000;
		b = 32'b00100111000001011011001011110111;
		correct = 32'b10110010000101101011010000010110;
		#400 //-4727752.0 * 1.8554475e-15 = -8.772096e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110101100100001001110000110010;
		b = 32'b00100010000100010101101101110110;
		correct = 32'b01011000001001000011100001000101;
		#400 //3.6663026e+32 * 1.9699583e-18 = 722246300000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010001101011110100001000111101;
		b = 32'b00100010110010110111011000110111;
		correct = 32'b00110101000010110100101001110101;
		#400 //94091320000.0 * 5.5148425e-18 = 5.1889884e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010000010110010011000110000010;
		b = 32'b01011010111001000011100011001100;
		correct = 32'b10101011110000011010000001001000;
		#400 //-4.2833844e-29 * 3.2119372e+16 = -1.3757962e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001001111110110001111001000000;
		b = 32'b01100010100101001000000111001001;
		correct = 32'b11101101000100011010110011001100;
		#400 //-2057160.0 * 1.369735e+21 = -2.817764e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111011010011000010001001001000;
		b = 32'b01011100110101100111011100001000;
		correct = 32'b11011000101010110000001110010011;
		#400 //-0.0031148363 * 4.8293217e+17 = -1504254700000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101000100010110111110001000100;
		b = 32'b00110000110110011110000001000000;
		correct = 32'b01011001111011010110110100001010;
		#400 //5.26961e+24 * 1.5852564e-09 = 8353682400000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000011111101100011110010000110;
		b = 32'b01101010010101111001101011100101;
		correct = 32'b10101110110011110110000111010001;
		#400 //-1.4472476e-36 * 6.516263e+25 = -9.430646e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001011111000111000110011010100;
		b = 32'b01110011111000011111010100011111;
		correct = 32'b01000000010010001101100010101000;
		#400 //8.7649114e-32 * 3.5804396e+31 = 3.1382236
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100010011001101010110000001111;
		b = 32'b01111100101001110100101010111011;
		correct = 32'b11011111100101101011110110010100;
		#400 //-3.12619e-18 * 6.949034e+36 = -2.1724001e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011111010001010010110111111100;
		b = 32'b00111001001011111000110111101010;
		correct = 32'b10011001000001110011011110111110;
		#400 //-4.175441e-20 * 0.00016742168 = -6.9905935e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100000011001110010011111000100;
		b = 32'b00000000111101110100110110100101;
		correct = 32'b10100001110111110100110101111010;
		#400 //-6.662599e+19 * 2.2711221e-38 = -1.5131576e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111100001010101101111001100101;
		b = 32'b10001010101000010101000011101100;
		correct = 32'b10000111010101110101011111000001;
		#400 //0.010429 * -1.5534175e-32 = -1.6200591e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001111011000011001010000101001;
		b = 32'b01010100100010100010111101101101;
		correct = 32'b10100100011100111000011101010001;
		#400 //-1.1121891e-29 * 4748009300000.0 = -5.2806843e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110101110000000001010011110101;
		b = 32'b10000111011111000010011111001010;
		correct = 32'b10111101101111010011001001111100;
		#400 //4.8698538e+32 * -1.8970066e-34 = -0.09238145
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101011011111010010010001000101;
		b = 32'b00111010111001111111011110101101;
		correct = 32'b11100110111001010110000010100011;
		#400 //-3.0602951e+26 * 0.0017697715 = -5.4160228e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000111110100010110001111101;
		b = 32'b11110111010111011001000100001000;
		correct = 32'b01101000110110001000011000100011;
		#400 //-1.8202538e-09 * -4.493903e+33 = 8.1800444e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101011110010110111100010100010;
		b = 32'b01010001001010001111000110011111;
		correct = 32'b00111101100001100100011100110101;
		#400 //1.44575e-12 * 45350515000.0 = 0.065565504
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110111011000111111111001011;
		b = 32'b11101110010110100001001101001000;
		correct = 32'b11101101110010010111011010100011;
		#400 //0.46191248 * -1.687276e+28 = -7.793739e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111000010000101101100010010110;
		b = 32'b10001110001111000110111000110101;
		correct = 32'b01000111000011110110101011110000;
		#400 //-1.5807789e+34 * -2.3225852e-30 = 36714.938
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110100010101111101110111100000;
		b = 32'b10100100101110000100000111000101;
		correct = 32'b11011001100110110101111011101110;
		#400 //6.841089e+31 * -7.99087e-17 = -5466624700000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000011010000101101010011000111;
		b = 32'b00001100010111011100100001011001;
		correct = 32'b00010000001010001100101000101010;
		#400 //194.83116 * 1.7085511e-31 = 3.32879e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001111010110111101001111110001;
		b = 32'b11101100100100011101011100001110;
		correct = 32'b00111100011110100111011101101101;
		#400 //-1.0838352e-29 * -1.4104785e+27 = 0.015287262
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111000010101001110101100110111;
		b = 32'b10001010110000110000100001000000;
		correct = 32'b00000011101000100011011000000111;
		#400 //-5.07638e-05 * -1.878092e-32 = 9.533908e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101110010010110010001010000100;
		b = 32'b11000000000011101010100100111111;
		correct = 32'b00101110111000100110011011100010;
		#400 //-4.6187512e-11 * -2.22908 = 1.0295566e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010010111001010111110010001111;
		b = 32'b01010010111111110111111110100110;
		correct = 32'b10100110011001010000100110000000;
		#400 //-1.4482638e-27 * 548679120000.0 = -7.946321e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010100000111110011100101000110;
		b = 32'b10100010001010110100100010010100;
		correct = 32'b10110110110101010001000011001100;
		#400 //2735442800000.0 * -2.3213244e-18 = -6.34985e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011100000110110111110010110011;
		b = 32'b01011001011000110001111001011111;
		correct = 32'b10110110000010011111001000000101;
		#400 //-5.144637e-22 * 3995513300000000.0 = -2.0555465e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111100101011000000001101001110;
		b = 32'b10001100011111000001000100111011;
		correct = 32'b11001001101010010101111011010101;
		#400 //7.145137e+36 * -1.9418559e-31 = -1387482.6
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001100111010111101110000011100;
		b = 32'b00011010000000100010110100001100;
		correct = 32'b00100111011011111101111010001110;
		#400 //123658460.0 * 2.691976e-23 = 3.328856e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110101011100110011000101010101;
		b = 32'b10111010001101111100001011000101;
		correct = 32'b01110000001011101001000101001010;
		#400 //-3.0828338e+32 * -0.0007009919 = 2.1610414e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010000000010010110011000101011;
		b = 32'b11101000101110011101001001011001;
		correct = 32'b10111001010001110111011101110101;
		#400 //2.7097193e-29 * -7.020144e+24 = -0.0001902262
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100111111101011001110001011;
		b = 32'b11100000100010000010101111110110;
		correct = 32'b11100110000001110111101100011111;
		#400 //2037.6107 * -7.849765e+19 = -1.5994766e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001111101111110010010001000011;
		b = 32'b11011110001001101101000001001010;
		correct = 32'b01101110011110010001101000010000;
		#400 //-6413649400.0 * -3.0050472e+18 = 1.9273319e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001010010001111001011100000010;
		b = 32'b01101011011110000100110111000011;
		correct = 32'b01110110010000011001011011101010;
		#400 //3270080.5 * 3.0018082e+26 = 9.816154e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101100011111000011101010101010;
		b = 32'b11111010011001000001011101111111;
		correct = 32'b01100111011000001011101101100110;
		#400 //-3.584392e-12 * -2.9608006e+35 = 1.061267e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101110010110000010010001110011;
		b = 32'b11000000110100110011111000110011;
		correct = 32'b00101111101100100101101010001111;
		#400 //-4.9145087e-11 * -6.6013427 = 3.2442357e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011010110110010011011101110010;
		b = 32'b11100011001110111110010010011010;
		correct = 32'b11111110100111110110110101111000;
		#400 //3.0570516e+16 * -3.4660136e+21 = -1.0595782e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111001111011110011000110000010;
		b = 32'b11001100111111101001101000000011;
		correct = 32'b01000111011011011110001100000110;
		#400 //-0.00045622519 * -133484570.0 = 60899.023
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011010001011110101111100011011;
		b = 32'b10110101110000011000000101101110;
		correct = 32'b01010000100001001000111101011110;
		#400 //-1.2340673e+16 * -1.441729e-06 = 17791906000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111100010101011110011110000111;
		b = 32'b00101000001000110111001101011001;
		correct = 32'b00100101000010001001001011001100;
		#400 //0.013055689 * 9.07333e-15 = 1.1845856e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100110010101111110001110111100;
		b = 32'b01000110110010011101010010011110;
		correct = 32'b10101101101010100011010100011100;
		#400 //-7.4901747e-16 * 25834.309 = -1.9350348e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010110000100001010100111110101;
		b = 32'b11001110010100101011100000000111;
		correct = 32'b10100100111011100010011011010010;
		#400 //1.1685856e-25 * -883818940.0 = -1.0328181e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010111100010010010100111010001;
		b = 32'b01100110101101101110001010010100;
		correct = 32'b00111110110000111111101001000010;
		#400 //8.863973e-25 * 4.3182516e+23 = 0.3827687
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010010010000100101110011101110;
		b = 32'b10010000100010000011001110110010;
		correct = 32'b00100011010011101101000100111100;
		#400 //-208695690000.0 * -5.372219e-29 = 1.12115895e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000111101100011101011101000;
		b = 32'b00011100100101000010011101100000;
		correct = 32'b10001110000011100111111111101101;
		#400 //-1.7915598e-09 * 9.803997e-22 = -1.7564445e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101001000001001100001111101111;
		b = 32'b01010101110111010000000101101010;
		correct = 32'b11111111011001010011101111000010;
		#400 //-1.0031467e+25 * 30374768000000.0 = -3.047035e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111010101110100000010010100;
		b = 32'b00111101000101111110100001111100;
		correct = 32'b01000100111111110111010100100100;
		#400 //55104.58 * 0.03708695 = 2043.6606
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011100101011001010011000000101;
		b = 32'b01100000000010011101111011111000;
		correct = 32'b11111101001110011111011001110000;
		#400 //-3.887699e+17 * 3.97386e+19 = -1.5449172e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111011010001111000010000011101;
		b = 32'b11111101001110110001110010001001;
		correct = 32'b11111001000100011101001110111110;
		#400 //0.0030443736 * -1.5544612e+37 = -4.7323605e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101101110111001011001101010010;
		b = 32'b00010110001101111011101010101001;
		correct = 32'b00000100100111100110010100011100;
		#400 //2.5090739e-11 * 1.4841522e-25 = 3.7238476e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111101111110110111000110100111;
		b = 32'b10110110000000011101111010111000;
		correct = 32'b00110100011111110001111000001101;
		#400 //-0.12277537 * -1.9352137e-06 = 2.3759658e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110010000100110100101101011101;
		b = 32'b10110110011110011111010110111101;
		correct = 32'b10101001000011111101000110110001;
		#400 //8.573662e-09 * -3.724693e-06 = -3.1934257e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110010010100101000010000100111;
		b = 32'b00001000111001101010100010000101;
		correct = 32'b00111011101111011010110101001111;
		#400 //4.1697033e+30 * 1.388224e-33 = 0.0057884823
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111100000000111100111000100010;
		b = 32'b01110101001010111100110000111111;
		correct = 32'b01110001101100001110011110110011;
		#400 //0.008044751 * 2.1777963e+32 = 1.751983e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001101001010101111000000111101;
		b = 32'b01001010011010010000111100001111;
		correct = 32'b00011000000110111001111010110110;
		#400 //5.267447e-31 * 3818435.8 = 2.0113409e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111000000011010001011001110010;
		b = 32'b10111011000101010110111100000011;
		correct = 32'b11110011101001001011011001111101;
		#400 //1.1446392e+34 * -0.0022801764 = -2.6099792e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000101001010000110001011100010;
		b = 32'b01001110101001101011111010111111;
		correct = 32'b11010100010110110101101100101011;
		#400 //-2694.1802 * 1398759300.0 = -3768509500000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110100001110011111001100100110;
		b = 32'b10110111000110100101001111101111;
		correct = 32'b01101011111000000011001001111001;
		#400 //-5.8929843e+31 * -9.198658e-06 = 5.4207547e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100001100010100000010100100111;
		b = 32'b00011010010011111000001111101010;
		correct = 32'b10111100010111111100001010010011;
		#400 //-3.1825274e+20 * 4.2913156e-23 = -0.01365723
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001001101000001001001000101011;
		b = 32'b00101101011010011001000100011001;
		correct = 32'b10110111100100101000000000001100;
		#400 //-1315397.4 * 1.3276735e-11 = -1.7464183e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110001111110110001000110111110;
		b = 32'b01110111111111010110111100110111;
		correct = 32'b01101010011110001000110110011011;
		#400 //7.3070785e-09 * 1.0280522e+34 = 7.512058e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011100111010110101101111000000;
		b = 32'b01001010110000001001100010010010;
		correct = 32'b01101000001100010001000100010101;
		#400 //5.2998e+17 * 6310985.0 = 3.344696e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110010001001111010011000111111;
		b = 32'b11000111010010011100111101100100;
		correct = 32'b01111010000001000010100101011000;
		#400 //-3.3206385e+30 * -51663.39 = 1.7155543e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010101011000110001011011011001;
		b = 32'b01101100111100010000010110110001;
		correct = 32'b11000010110101011100110110001111;
		#400 //-4.586031e-26 * 2.331024e+27 = -106.90148
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110010000100100010011011101001;
		b = 32'b10011101001010110000011000011101;
		correct = 32'b01001111110000110100011011110110;
		#400 //-2.8948385e+30 * -2.2634822e-21 = 6552415000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101000110111011011010011100000;
		b = 32'b10110110001011101010111110010011;
		correct = 32'b10011111100101110100100011111110;
		#400 //2.4614371e-14 * -2.6030218e-06 = -6.407174e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000110000010011110011010010000;
		b = 32'b11000011011111110100010000001110;
		correct = 32'b11001010000010011000000101010010;
		#400 //8825.641 * -255.26584 = -2252884.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101100101000011010110001001100;
		b = 32'b10111000010101101111110001001001;
		correct = 32'b10100101100001111100010101011011;
		#400 //4.595024e-12 * -5.1256535e-05 = -2.35525e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001111101011001101011010100100;
		b = 32'b11000010101000101111001110001010;
		correct = 32'b01010010110111000000100010000001;
		#400 //-5799495700.0 * -81.47566 = 472517740000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010010010011111111010000011100;
		b = 32'b01111011100010000110100100001111;
		correct = 32'b01001110010111011001111000001100;
		#400 //6.561857e-28 * 1.4165664e+36 = 929530600.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000011011110010110111011111010;
		b = 32'b01001110111111010101101101011111;
		correct = 32'b11010010111101101101101110110100;
		#400 //-249.4335 * 2125311900.0 = -530123980000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010100000100110011110000100111;
		b = 32'b11011101110000101111010011010000;
		correct = 32'b01110010011000000100000011000101;
		#400 //-2529477500000.0 * -1.7560102e+18 = 4.4417884e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101010001101001000000010011110;
		b = 32'b10011011101110010111101100100101;
		correct = 32'b10000110100000101100011111000110;
		#400 //1.6031835e-13 * -3.0685263e-22 = -4.9194106e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101101110000100001000111011100;
		b = 32'b00011111000010011110011100111000;
		correct = 32'b10001101010100010001010110101111;
		#400 //-2.2063178e-11 * 2.9202138e-20 = -6.44292e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001111101111110111010011101011;
		b = 32'b00110001101111101111010010011101;
		correct = 32'b10000010000011101100111110110111;
		#400 //-1.887909e-29 * 5.557537e-09 = -1.0492124e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000010010110011111001010011111;
		b = 32'b11000011010101000001100010110100;
		correct = 32'b11000110001101001001000111110100;
		#400 //54.486935 * -212.0965 = -11556.488
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001010111110001011110111001111;
		b = 32'b00001110100010100101000100010100;
		correct = 32'b00011010000001100110010100011001;
		#400 //8150759.5 * 3.4097702e-30 = 2.7792217e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110010110111111101001000000011;
		b = 32'b01110001011010000101110110111101;
		correct = 32'b01100100110010110010100001000111;
		#400 //2.6056119e-08 * 1.1506215e+30 = 2.998073e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100110101111010011001010100;
		b = 32'b00111001000100000011100101111101;
		correct = 32'b00111110011100101111101111111001;
		#400 //1725.1978 * 0.00013754326 = 0.23728932
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010100010001100000010110101110;
		b = 32'b10111110010100100110111010001010;
		correct = 32'b10010011001000101100011000101010;
		#400 //9.9975655e-27 * -0.2054998 = -2.0544977e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100101011010010001100100010101;
		b = 32'b11110111110001100101100101000010;
		correct = 32'b01011101101101001001101010101100;
		#400 //-2.0218027e-16 * -8.0459777e+33 = 1.6267379e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101101100001011000111110010011;
		b = 32'b01100010100010100000111100110001;
		correct = 32'b01010000100100000000111010100100;
		#400 //1.518411e-11 * 1.2733727e+21 = 19335029000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100000111000011100100100111001;
		b = 32'b00101111000101100001110110110110;
		correct = 32'b01010000100001000110011000011100;
		#400 //1.3015678e+20 * 1.3652976e-10 = 17770275000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100011000001110011100100001001;
		b = 32'b01001100110101000011000101101101;
		correct = 32'b00110000011000000010101010101110;
		#400 //7.330442e-18 * 111250280.0 = 8.1551377e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101110001101110101101000001111;
		b = 32'b10111111100011100001010011001110;
		correct = 32'b11101110010010111000010110110110;
		#400 //1.4186158e+28 * -1.1100099 = -1.5746776e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001101100111111100111010100110;
		b = 32'b11011101000011100011101101000001;
		correct = 32'b11101011001100011001001100111011;
		#400 //335140030.0 * -6.4055355e+17 = -2.1467515e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001010011111111100110111110101;
		b = 32'b01010010101110001011111111011011;
		correct = 32'b00011101101110001001101110111110;
		#400 //1.23165396e-32 * 396746400000.0 = 4.886543e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001101010111011111000001001011;
		b = 32'b10110110100010010110001000001010;
		correct = 32'b01000100011011100011010100101110;
		#400 //-232719540.0 * -4.0943314e-06 = 952.83093
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101101001101000000111010010100;
		b = 32'b01000000000000010000000101100001;
		correct = 32'b11101101101101010111100010100010;
		#400 //-3.482808e+27 * 2.0157092 = -7.020328e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100000111101001111001011000100;
		b = 32'b00110110100011110111011000100000;
		correct = 32'b10011000000010010100010010100010;
		#400 //-4.1495857e-19 * 4.2754837e-06 = -1.7741486e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000010001010001001000011100100;
		b = 32'b11010011011010000010101000000000;
		correct = 32'b00010110000110001101111011110110;
		#400 //-1.2384272e-37 * -997137060000.0 = 1.2348816e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111011100010101010100111001000;
		b = 32'b00011000100100000110000100110111;
		correct = 32'b00010100100111000110100001010001;
		#400 //0.0042316653 * 3.732129e-24 = 1.579312e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110011000111000111100010011010;
		b = 32'b01010110111010010011110001110000;
		correct = 32'b01001010100011101000111010110101;
		#400 //3.6431267e-08 * 128222890000000.0 = 4671322.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100001010011000101010000001101;
		b = 32'b01001000011110111111011001111100;
		correct = 32'b10101010010010010001101100100100;
		#400 //-6.922913e-19 * 258009.94 = -1.7861803e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100011010000001100111000010101;
		b = 32'b00111100010101001001101001101000;
		correct = 32'b11100000001000000001111011110100;
		#400 //-3.5566246e+21 * 0.012976266 = -4.615171e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111000011111111010011001110000;
		b = 32'b10110010011000111110111001111100;
		correct = 32'b10101011011000111001111010111110;
		#400 //6.0951745e-05 * -1.3267364e-08 = -8.08669e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101110001011111100010110101010;
		b = 32'b00100011000101001011000101011010;
		correct = 32'b11010001110011000011000000010111;
		#400 //-1.359971e+28 * 8.060652e-18 = -109622520000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101110010001000110111010010100;
		b = 32'b11110100011101111011011001001000;
		correct = 32'b01100011001111100001001010001111;
		#400 //-4.4663453e-11 * -7.850308e+31 = 3.5062187e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101000111010001001100011100010;
		b = 32'b00011000101111100001001000111000;
		correct = 32'b11000010001011001011001000000101;
		#400 //-8.787274e+24 * 4.9132245e-24 = -43.173847
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010010111111101001011010110101;
		b = 32'b11101010011110110101111100001010;
		correct = 32'b10111101111110011111110001000111;
		#400 //1.6066806e-27 * -7.5972298e+25 = -0.12206321
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111100001100010000100101100110;
		b = 32'b10110010100011010111000110101010;
		correct = 32'b01101111010000111010000110010000;
		#400 //-3.6769087e+36 * -1.6466249e-08 = 6.0544894e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101010000101101011100011010011;
		b = 32'b10000011111100000110000110100010;
		correct = 32'b00101110100011011000011011000001;
		#400 //-4.555292e+25 * -1.4128348e-36 = 6.435875e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011100100111110010111000001111;
		b = 32'b10110011110010011111010101100000;
		correct = 32'b10010000111110110010011101111001;
		#400 //1.0533643e-21 * -9.404425e-08 = -9.906286e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110110011111000100010110100000;
		b = 32'b00010110101001101101001111011011;
		correct = 32'b01001101101001000110010111101011;
		#400 //1.2791709e+33 * 2.6952446e-25 = 344767840.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001010000011110011101111110100;
		b = 32'b11000000100010110000100011010000;
		correct = 32'b11001011000110111001010011110111;
		#400 //2346749.0 * -4.3448257 = -10196215.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100100101101101011100000100111;
		b = 32'b11000001001010110011001110101101;
		correct = 32'b11100110011101000110001111001000;
		#400 //2.6964616e+22 * -10.700116 = -2.8852452e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010010111011110001111110000001;
		b = 32'b01000001111000111101001110100110;
		correct = 32'b11010101010101001100111010100001;
		#400 //-513512870000.0 * 28.478344 = -14623996000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101111100000001100111101001111;
		b = 32'b11010101110100100000001110110101;
		correct = 32'b11000101110100110101011111011001;
		#400 //2.3430366e-10 * -28864170000000.0 = -6762.981
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011111000111111101000101001010;
		b = 32'b00101010100010001010111110010111;
		correct = 32'b10001010001010101010100110011011;
		#400 //-3.384268e-20 * 2.4280293e-13 = -8.2171015e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101110101111000101111110000011;
		b = 32'b01001101111110001001110110110000;
		correct = 32'b01111101001101101111000010001111;
		#400 //2.9149324e+28 * 521385470.0 = 1.5198034e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011001100101010110010111010101;
		b = 32'b10100101001000110100110000100101;
		correct = 32'b00111111001111101001100010001101;
		#400 //-5256467000000000.0 * -1.4163795e-16 = 0.74451524
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001110101100100011101001111001;
		b = 32'b11110011100001111010010110101010;
		correct = 32'b11000010101111001110000001011000;
		#400 //4.3936695e-30 * -2.1494145e+31 = -94.43817
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011011111011010000101011110100;
		b = 32'b10101001010100100010000110000101;
		correct = 32'b00000101110000101001001000000110;
		#400 //-3.921544e-22 * -4.665844e-14 = 1.8297313e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111010100011111000010101011101;
		b = 32'b10000110000111111110001100100010;
		correct = 32'b10000001001100110100011001010110;
		#400 //0.001094978 * -3.0071447e-35 = -3.292757e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011000011001110000100100011010;
		b = 32'b10010100010011100010110011011001;
		correct = 32'b00101101001110100001000111001100;
		#400 //-1016105100000000.0 * -1.0409187e-26 = 1.0576828e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011100111100001010100011101101;
		b = 32'b00111000110000110011110010111111;
		correct = 32'b01010110001101111000100111001000;
		#400 //5.4191784e+17 * 9.3096394e-05 = 50450600000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010111101101000010010011110110;
		b = 32'b01111100000111111010100000010001;
		correct = 32'b11010100011000001011001001110010;
		#400 //-1.1641558e-24 * 3.315936e+36 = -3860266000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111110111101000110011001101100;
		b = 32'b00010011100110100100101110001110;
		correct = 32'b10010011000100110100110110111111;
		#400 //-0.47734392 * 3.894957e-27 = -1.859234e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111000011011001111110110000;
		b = 32'b01000111000010100100110000010110;
		correct = 32'b01001110100110010000010001011001;
		#400 //36255.688 * 35404.086 = 1283599500.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100011111100111100111111110001;
		b = 32'b10010110111011110101101101001010;
		correct = 32'b10111011011000111111011000010011;
		#400 //8.995085e+21 * -3.8670144e-25 = -0.0034784123
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100010100101101110100011101000;
		b = 32'b11011011111000111001110011001111;
		correct = 32'b10111111000001100010110011110110;
		#400 //4.090418e-18 * -1.28134465e+17 = -0.52412355
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000101001011100011010011101100;
		b = 32'b01101010100011000001100001101110;
		correct = 32'b10110000001111101010101100100010;
		#400 //-8.191161e-36 * 8.468249e+25 = -6.936479e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111111010010100001001001000010;
		b = 32'b10110101000101100110011100001010;
		correct = 32'b01110100111011010111000000010000;
		#400 //-2.6859886e+38 * -5.6029296e-07 = 1.5049405e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011000100000101100001100000001;
		b = 32'b10001000010111100001111011111100;
		correct = 32'b10100001011000101110100111011101;
		#400 //1150192400000000.0 * -6.6842117e-34 = -7.6881294e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010000011000010011010110111110;
		b = 32'b11011110101100101100010101010001;
		correct = 32'b10101111100111010100010011110100;
		#400 //4.4414827e-29 * -6.4408957e+18 = -2.8607128e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011101011111110110100110001111;
		b = 32'b01100011001111011110000111100011;
		correct = 32'b01000001001111010111001001001101;
		#400 //3.3803542e-21 * 3.5027115e+21 = 11.840405
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101010011101000101110111111111;
		b = 32'b01010010000011011011111010111111;
		correct = 32'b00111101000001110100110111011010;
		#400 //2.1704165e-13 * 152197640000.0 = 0.03303323
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001111101000011110101010001000;
		b = 32'b00010010100001001101010010111100;
		correct = 32'b00100010101010000000011011110111;
		#400 //5433004000.0 * 8.382814e-28 = 4.5543866e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011100001100111010111101011101;
		b = 32'b11110001000001100011010100111100;
		correct = 32'b01001101101111000110011001010000;
		#400 //-5.9452784e-22 * -6.645656e+29 = 395102720.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110001111000011011100101111011;
		b = 32'b01000011100110001100000110111000;
		correct = 32'b11110110000001101011000011110000;
		#400 //-2.2354675e+30 * 305.51343 = -6.829653e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010100101100011000010001110101;
		b = 32'b01000100000100010101101011110001;
		correct = 32'b01011001010010011001011000101100;
		#400 //6099452000000.0 * 581.42096 = 3546349000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000101001001110100110111010010;
		b = 32'b11010110110011001100010000010111;
		correct = 32'b10011100100001011101001000101010;
		#400 //7.8665956e-36 * -112571286000000.0 = -8.855528e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010111000000100001001100110011;
		b = 32'b00101010011000111110101011101001;
		correct = 32'b11000001111001111001110011000100;
		#400 //-143018970000000.0 * 2.0243151e-13 = -28.951546
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000101000010010011101110111011;
		b = 32'b11001011001011111001011110001101;
		correct = 32'b01010000101111000100001000100101;
		#400 //-2195.7332 * -11507597.0 = 25267612000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000100011010010100000011001100;
		b = 32'b01110111011101100001001001001110;
		correct = 32'b10111100011000000011010011110010;
		#400 //-2.7418772e-36 * 4.990923e+33 = -0.013684498
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100100110110111101110001111000;
		b = 32'b01010110001011011001110000110001;
		correct = 32'b01111011100101010001101000100010;
		#400 //3.2445787e+22 * 47721587000000.0 = 1.5483645e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001010111110100000101001011101;
		b = 32'b00010001000001000101010011010110;
		correct = 32'b10011100100000010100000000110100;
		#400 //-8193326.5 * 1.0439106e-28 = -8.5531e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000111001111001110100011100000;
		b = 32'b11111000101000100101100001101111;
		correct = 32'b01000000011011111001100100111111;
		#400 //-1.4211984e-34 * -2.6342054e+34 = 3.7437284
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111000001001011100010110000011;
		b = 32'b10110001001011101001010111111001;
		correct = 32'b01101001111000100001101010111000;
		#400 //-1.3448984e+34 * -2.5405582e-09 = 3.4167926e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001101010000110001000111011100;
		b = 32'b00111101010110010111011010101010;
		correct = 32'b10001011001001011011010010001111;
		#400 //-6.011051e-31 * 0.053091682 = -3.191368e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001000101100111010101110011000;
		b = 32'b01011111101000110010010111011101;
		correct = 32'b00101000111001010000000110101001;
		#400 //1.0813512e-33 * 2.351209e+19 = 2.5424827e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001000101001001110011001000001;
		b = 32'b00111011101111101111100001010011;
		correct = 32'b11000100111101100000010110110010;
		#400 //-337714.03 * 0.0058279424 = -1968.178
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100011101001000010111001000010;
		b = 32'b11101000111010100001111011111101;
		correct = 32'b01001101000101100010011000101000;
		#400 //-1.7800507e-17 * -8.844843e+24 = 157442690.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000110000101001100110000110101;
		b = 32'b11100011000001001011010111100000;
		correct = 32'b10101001100110100100011000000100;
		#400 //2.7985734e-35 * -2.4480757e+21 = -6.8511196e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101110110100111110110101110110;
		b = 32'b00101111010110100101001001101011;
		correct = 32'b10011110101101001011110001110001;
		#400 //-9.6373506e-11 * 1.9856265e-10 = -1.9136179e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011101100111001001010000111110;
		b = 32'b00111111011000100110010010001000;
		correct = 32'b11011101100010100111100001011100;
		#400 //-1.4103389e+18 * 0.8843465 = -1.2472283e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110101111111010111010001001101;
		b = 32'b00101110101100001000110111010001;
		correct = 32'b00100101001011101100110001011101;
		#400 //1.8883817e-06 * 8.028745e-11 = 1.5161335e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011000010101011111111011100101;
		b = 32'b01010101011100010001000101000000;
		correct = 32'b00101110010010011000001101100001;
		#400 //2.7658294e-24 * 16566024000000.0 = 4.5818797e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001000010010101101011011100011;
		b = 32'b11000111010010010000111000101111;
		correct = 32'b01010000000111110100110111110101;
		#400 //-207707.55 * -51470.184 = 10690745000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101101000011110000011101110010;
		b = 32'b01000100100010111000101101001110;
		correct = 32'b10110010000110111110110110111111;
		#400 //-8.130262e-12 * 1116.3533 = -9.076245e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000101011110010110100011110110;
		b = 32'b11110001110000110011101000111011;
		correct = 32'b11110111101111100011001110101111;
		#400 //3990.56 * -1.9334391e+30 = -7.715505e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011100011000110011101011001111;
		b = 32'b01001000100100011010100010110110;
		correct = 32'b11100101100000010100101000001111;
		#400 //-2.5583792e+17 * 298309.7 = -7.631893e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000101010111111011010110001011;
		b = 32'b11110100000111000011101001000010;
		correct = 32'b01111010000010001000010110001010;
		#400 //-3579.3464 * -4.9510493e+31 = 1.7721522e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011011000100000001100111000101;
		b = 32'b01011000011110101001000110100010;
		correct = 32'b11110100000011010000101100100100;
		#400 //-4.056073e+16 * 1102013600000000.0 = -4.4698475e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111100011001001111001010001010;
		b = 32'b11100101001001010011011010111100;
		correct = 32'b11100010000100111100000101000110;
		#400 //0.013973841 * -4.876251e+22 = -6.8139955e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010110000000110100110001010001;
		b = 32'b11100110011000001100011101101100;
		correct = 32'b00111100111001101001001000011101;
		#400 //-1.0606177e-25 * -2.653722e+23 = 0.028145844
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100010110001111101000010110000;
		b = 32'b10110110000010110100000110001111;
		correct = 32'b01011001010110010110001011110110;
		#400 //-1.8429698e+21 * -2.0750774e-06 = 3824305000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000101011010111001100000100110;
		b = 32'b11110010010011011110100010111101;
		correct = 32'b01111000001111010111111100000110;
		#400 //-3769.5093 * -4.0784506e+30 = 1.5373757e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010100001100111110000100101110;
		b = 32'b00111110011001101111100110110011;
		correct = 32'b00010011001000100100101111000011;
		#400 //9.0815994e-27 * 0.2255619 = 2.0484628e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011010110101111110101000010010;
		b = 32'b11100110001011110110010000111110;
		correct = 32'b11000001100100111110110110001110;
		#400 //8.9300077e-23 * -2.0706582e+23 = -18.490993
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010000111111110010101010001110;
		b = 32'b01111111010100111100101101101111;
		correct = 32'b11010000110100110001101011011000;
		#400 //-1.0064533e-28 * 2.815234e+38 = -28334014000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110000110000010000111101111010;
		b = 32'b10110001000101001110011011010000;
		correct = 32'b01100010011000001001011000000111;
		#400 //-4.7799454e+29 * -2.1668036e-09 = 1.0357203e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001111110000110101000001001101;
		b = 32'b11101100111011000100110111101000;
		correct = 32'b10111101001101000100100101110111;
		#400 //1.9259415e-29 * -2.2853952e+27 = -0.044015374
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111001010110000010111010101110;
		b = 32'b01100001101101100101011110100011;
		correct = 32'b01011011100110011111101100110001;
		#400 //0.00020616755 * 4.204528e+20 = 8.668372e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111110000011011000101011010000;
		b = 32'b10111010101100110110001010101101;
		correct = 32'b00111001010001100101110100111100;
		#400 //-0.13822484 * -0.0013686024 = 0.00018917484
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001110000111010101111100000111;
		b = 32'b10100010100101111111100000110111;
		correct = 32'b00110001001110101101011101000110;
		#400 //-660062660.0 * -4.119144e-18 = 2.718893e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111010101101101101001000110;
		b = 32'b01110001001010010101011011111101;
		correct = 32'b01111001000011100001111100011010;
		#400 //55002.273 * 8.385301e+29 = 4.612106e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101110101011110111001101001011;
		b = 32'b01001010010101001011010010010011;
		correct = 32'b01111001100100011100011100111100;
		#400 //2.7149629e+28 * 3484964.8 = 9.46155e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110101001111110110011011100000;
		b = 32'b10011110000010010001101110110111;
		correct = 32'b11010011110011010000010110001101;
		#400 //2.4263068e+32 * -7.258451e-21 = -1761122800000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000000101110011101100000111111;
		b = 32'b00110000101100110011000000111101;
		correct = 32'b10110010000000100001010100111001;
		#400 //-5.807647 * 1.3037674e-09 = -7.571821e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111100101011101011010111001110;
		b = 32'b01010111000111101011101001111001;
		correct = 32'b11010100010110001010011011110000;
		#400 //-0.021326926 * 174523730000000.0 = -3722054700000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111100001010000111101101000010;
		b = 32'b10001110010010100110100010000110;
		correct = 32'b10001011000001010011011000001100;
		#400 //0.010283293 * -2.4948749e-30 = -2.565553e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110101011000001001000010000010;
		b = 32'b00101001000100001000110100100001;
		correct = 32'b11011110111111011001101000101011;
		#400 //-2.846693e+32 * 3.2096833e-14 = -9.136983e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110111010100111000010100001110;
		b = 32'b11010111111110011000000100001100;
		correct = 32'b11001111110011100010011100001011;
		#400 //1.2607559e-05 * -548665300000000.0 = -6917330400.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010010111010000110010010100011;
		b = 32'b01011001010101111101000110110110;
		correct = 32'b10101100110000111110101011100100;
		#400 //-1.4666067e-27 * 3796731200000000.0 = -5.5683114e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011010110101101110001100110101;
		b = 32'b01101011011111010111110110010111;
		correct = 32'b11000110110101001100011111110111;
		#400 //-8.88754e-23 * 3.0645131e+26 = -27235.982
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000011001010010101010100010111;
		b = 32'b11011110110100111101011100101101;
		correct = 32'b00100010100011000001111101110110;
		#400 //-4.9762315e-37 * -7.6323595e+18 = 3.7980387e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010101010100011010100011100001;
		b = 32'b00101110110000101010011110001011;
		correct = 32'b11000100100111110110101100110010;
		#400 //-14407704000000.0 * 8.85186e-11 = -1275.3499
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001100110000110110110111111010;
		b = 32'b00100011101011011101010011000100;
		correct = 32'b00110001000001001011001110111111;
		#400 //102461390.0 * 1.8846807e-17 = 1.9310702e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010111000011011101111110000111;
		b = 32'b10001001011011010110111010001011;
		correct = 32'b00100001000000111001010100110011;
		#400 //-155991180000000.0 * -2.8579814e-33 = 4.458199e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111111101011101111111001011101;
		b = 32'b11010011001000001010110100100001;
		correct = 32'b11010011010110111010101010100101;
		#400 //1.3671376 * -690099400000.0 = -943460800000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011001110111011100100001110100;
		b = 32'b00000110011001000111101011011000;
		correct = 32'b00100000110001011111000011110100;
		#400 //7803296300000000.0 * 4.2972285e-35 = 3.3532548e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100010110111110000100010001110;
		b = 32'b11010101011101100001110000101001;
		correct = 32'b10111000110101100110101011000001;
		#400 //6.045333e-18 * -16912550000000.0 = -0.000102242
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011110010001000000101010001110;
		b = 32'b10100100001011110011100000101101;
		correct = 32'b00000011000001100010111000111100;
		#400 //-1.0378336e-20 * -3.799466e-17 = 3.9432135e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100100011110110101101110010010;
		b = 32'b01110111100011110001011001110010;
		correct = 32'b01011100100011000111111000110000;
		#400 //5.4504512e-17 * 5.804326e+33 = 3.1636193e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000111000011000101011011001010;
		b = 32'b10101010011100011101111100110110;
		correct = 32'b00110010000001001001100000010001;
		#400 //-35926.79 * -2.1482542e-13 = 7.717987e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111001010000000001101111100110;
		b = 32'b01011101110001011000010010011111;
		correct = 32'b11010111100101000011100011111110;
		#400 //-0.0001832094 * 1.7790844e+18 = -325945000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010111001111111110111001101111;
		b = 32'b10010101110111001110001111000101;
		correct = 32'b00101101101001011001101110101100;
		#400 //-211030790000000.0 * -8.921665e-26 = 1.882746e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110101111100000000010011100111;
		b = 32'b10111110010100110001111001111100;
		correct = 32'b10110100110001011111000010011111;
		#400 //1.788282e-06 * -0.20617098 = -3.6869184e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011101111001000111011000100001;
		b = 32'b11000000010001000100000011000011;
		correct = 32'b00011110101011110010010000111101;
		#400 //-6.047324e-21 * -3.0664527 = 1.8543834e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101100100101110001000001110011;
		b = 32'b11110101100000111110011011110100;
		correct = 32'b11100010100110111010101101100111;
		#400 //4.2935044e-12 * -3.344117e+32 = -1.4357981e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010110101110011111111010001110;
		b = 32'b11000110010101001110101100000101;
		correct = 32'b11011101100110101011000110001110;
		#400 //102251480000000.0 * -13626.755 = -1.3933558e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110111110111000010010100010000;
		b = 32'b10011011100101011100011001111010;
		correct = 32'b01010100000000001100110001000000;
		#400 //-8.930133e+33 * -2.4778245e-22 = 2212730200000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010101010011010101100101100111;
		b = 32'b11011001100001010100000011100010;
		correct = 32'b00101111010101011100011011111100;
		#400 //-4.1469946e-26 * -4688439000000000.0 = 1.944293e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011011010110110001100001010010;
		b = 32'b00101101001011100111000010010110;
		correct = 32'b11001001000101010100101011100011;
		#400 //-6.166976e+16 * 9.915754e-12 = -611502.2
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100000010100100011001111100110;
		b = 32'b11011000001101000000000011101011;
		correct = 32'b00111001000100111100110100111111;
		#400 //-1.7804864e-19 * -791664140000000.0 = 0.00014095473
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111000100010010001000001010101;
		b = 32'b00100110111100000011110101011010;
		correct = 32'b01100000000000001010000000101001;
		#400 //2.2239873e+34 * 1.6669975e-15 = 3.7073812e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001011110000001010110100011101;
		b = 32'b01011111001100011011110001010101;
		correct = 32'b00101011100001011100010101110000;
		#400 //7.421618e-32 * 1.2807205e+19 = 9.505018e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011000100001000010101111101111;
		b = 32'b11001001010010011101010000100010;
		correct = 32'b11100010010100000110100000001001;
		#400 //1162593800000000.0 * -826690.1 = -9.611048e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111000011100011011011010010111;
		b = 32'b11100110101110101100000010100000;
		correct = 32'b01011111101100000101010010001010;
		#400 //-5.7628928e-05 * -4.4095673e+23 = 2.5411864e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111101100001110100001111111110;
		b = 32'b01100011101111000010101100100100;
		correct = 32'b11100001110001101101100101110100;
		#400 //-0.06604765 * 6.942193e+21 = -4.5851556e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110110100100011100111111000001;
		b = 32'b01100110010010101101000111011010;
		correct = 32'b01011101011001110000101011101010;
		#400 //4.3455225e-06 * 2.3944728e+23 = 1.0405235e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110011010000110010010100101101;
		b = 32'b11000001001100001001101000111010;
		correct = 32'b10110101000001101001111100100000;
		#400 //4.5435787e-08 * -11.037653 = -5.015045e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110100011100010010000110011110;
		b = 32'b01100101010011010101111110001110;
		correct = 32'b01011010010000010111000111101101;
		#400 //2.2457104e-07 * 6.0615488e+22 = 1.3612483e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010111000000111100010000111110;
		b = 32'b11101101000011001011110001011110;
		correct = 32'b11000100100100001110000010001101;
		#400 //4.2576075e-25 * -2.7222265e+27 = -1159.0172
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010100001001101000011010001010;
		b = 32'b00110101111011100101100111101011;
		correct = 32'b11001010100110110000101110010010;
		#400 //-2860887000000.0 * 1.7758551e-06 = -5080521.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111101001111000101000010010101;
		b = 32'b00000101100010100010101100100001;
		correct = 32'b01000011010010110100011001010100;
		#400 //1.5644579e+37 * 1.29933e-35 = 203.27472
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001100000010100011101111010001;
		b = 32'b00100100110101010101011000101010;
		correct = 32'b10110001011001100110010010010111;
		#400 //-36237124.0 * 9.251999e-17 = -3.3526584e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000001010010010001110001101000;
		b = 32'b11110000010111011101001001001100;
		correct = 32'b00110010001011100100001010111011;
		#400 //-3.693825e-38 * -2.7460168e+29 = 1.0143306e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001010100001101110110001110100;
		b = 32'b01011111001110011110101011111001;
		correct = 32'b01101010010000111111100101101110;
		#400 //4421178.0 * 1.3396794e+19 = 5.922961e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010101010110000001010000111011;
		b = 32'b00001110110001001100101001100101;
		correct = 32'b00100100101001100001101001010010;
		#400 //14848838000000.0 * 4.851263e-30 = 7.203561e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001011011010001001010100111100;
		b = 32'b11011011000110011001110100101110;
		correct = 32'b10100111000010111000111111111110;
		#400 //4.4793846e-32 * -4.3238492e+16 = -1.9368183e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000110110100101111001101000001;
		b = 32'b01100111101110011100100101000011;
		correct = 32'b10101111000110010001011110100010;
		#400 //-7.935065e-35 * 1.7547008e+24 = -1.3923665e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011110100011011111000110101011;
		b = 32'b11111100101001110101011000000111;
		correct = 32'b11011011101110011001000010110011;
		#400 //1.5028907e-20 * -6.9508673e+36 = -1.0446394e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111001011000111110000111101101;
		b = 32'b11011010101000111101110000100001;
		correct = 32'b11010100100100011101110011001101;
		#400 //0.00021732571 * -2.3061228e+16 = -5011797400000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011010110000000011011001101111;
		b = 32'b10101010011101101111000111000100;
		correct = 32'b00000101101110010110100111010101;
		#400 //-7.949728e-23 * -2.1933068e-13 = 1.7436193e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000001000101100101001111110111;
		b = 32'b01011100100100010010100111100011;
		correct = 32'b00011110001010100111110001001111;
		#400 //2.761089e-38 * 3.268794e+17 = 9.0254315e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111100001001111110101111001001;
		b = 32'b11011100011000110101011100101001;
		correct = 32'b01011001000101010001111100111111;
		#400 //-0.010249087 * -2.5596261e+17 = 2623383000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101010100111110110001000000111;
		b = 32'b10100011111110000011111010000011;
		correct = 32'b11001111000110101000110111100010;
		#400 //9.634106e+25 * -2.6914689e-17 = -2592989700.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100110010001101000100111101100;
		b = 32'b00110100000101110111000111101000;
		correct = 32'b01011010111010101110011101100010;
		#400 //2.343932e+23 * 1.410441e-07 = 3.3059776e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001000001011100110110000110000;
		b = 32'b11100010001000010100100101011101;
		correct = 32'b10101010110110111100100000001101;
		#400 //5.2488394e-34 * -7.4380304e+20 = -3.9041028e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000000111101111100111110010011;
		b = 32'b01000111110000111001101001101011;
		correct = 32'b01001001001111010101100010010111;
		#400 //7.7440886 * 100148.836 = 775561.44
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110010011000110001001000111010;
		b = 32'b00010011000100011100001101010000;
		correct = 32'b11000110000000010100101010010001;
		#400 //-4.4976084e+30 * 1.839787e-27 = -8274.642
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111100111000010100001101110011;
		b = 32'b00111111000001001011101010001000;
		correct = 32'b11111100011010011001010111010100;
		#400 //-9.3570786e+36 * 0.51847124 = -4.8513762e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000011011111010111111110100;
		b = 32'b10011000000011001111110011000111;
		correct = 32'b00001001000001000000000011100101;
		#400 //-8.719774e-10 * -1.8222196e-24 = 1.5889343e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001101100110010000011011011100;
		b = 32'b00110100110001010010110111111111;
		correct = 32'b10000010111010111011101110001100;
		#400 //-9.431004e-31 * 3.6727576e-07 = -3.4637793e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100011001010111010111101010001;
		b = 32'b01111110100111110011011111010010;
		correct = 32'b01100010010101011000111010100110;
		#400 //9.307053e-18 * 1.0581854e+38 = 9.8485885e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010011011010100011110001110011;
		b = 32'b01001101111111001000100000111110;
		correct = 32'b00100001111001110001000000101010;
		#400 //2.9564756e-27 * 529598400.0 = 1.5657447e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000010101001111000111001010101;
		b = 32'b00011111100010111100010010000010;
		correct = 32'b00100010101101101111010111001100;
		#400 //83.77799 * 5.9193885e-20 = 4.9591446e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010100100010100001000100001110;
		b = 32'b00111111010000000101010110001010;
		correct = 32'b01010100010011110111010111011001;
		#400 //4743933000000.0 * 0.7513052 = 3564141500000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011100111111011001100011000;
		b = 32'b11000011000111101111001100111100;
		correct = 32'b01001111010001100101000010001010;
		#400 //-20932144.0 * -158.95013 = 3327167000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111011110010111010010000001;
		b = 32'b10111011010000111100110011100111;
		correct = 32'b11000011001111101100101101101000;
		#400 //63860.504 * -0.002987677 = -190.79456
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010011001111011101001001111011;
		b = 32'b10000100101010110010111001110000;
		correct = 32'b10011000011111011101110000001110;
		#400 //815280100000.0 * -4.0244553e-36 = -3.2810583e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101010011101111011110101010001;
		b = 32'b00100101110000110010011100011111;
		correct = 32'b01010000101111001101101100010001;
		#400 //7.4874675e+25 * 3.3853617e-16 = 25347787000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101011000011111100011000111101;
		b = 32'b10111111101000101110011101011101;
		correct = 32'b00101011001101101111101011000101;
		#400 //-5.1078916e-13 * -1.2726856 = 6.50074e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001010011010101010110001010111;
		b = 32'b01101011001111100010100101001010;
		correct = 32'b10110110001011100101000111000010;
		#400 //-1.1299104e-32 * 2.2989089e+26 = -2.597561e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101011100011101001100000100101;
		b = 32'b11000100111001010011111100100011;
		correct = 32'b01110000111111110110001010001000;
		#400 //-3.447719e+26 * -1833.973 = 6.3230236e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011111010100100100101001101010;
		b = 32'b11001001101011110000110011100111;
		correct = 32'b11101001100011111100101101111000;
		#400 //1.515304e+19 * -1434012.9 = -2.1729656e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111100000110001011111101110101;
		b = 32'b00001011100101001100100001101010;
		correct = 32'b10001000001100011000110010001001;
		#400 //-0.009322991 * 5.7309076e-32 = -5.34292e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101000000110100111011010011111;
		b = 32'b00011011001000011110010100100001;
		correct = 32'b00000011110000110101110110110100;
		#400 //8.574439e-15 * 1.3391643e-22 = 1.1482583e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011111100101110011111001101111;
		b = 32'b01100010010101011111101001011001;
		correct = 32'b11000010011111001101010110110100;
		#400 //-6.4054275e-20 * 9.86799e+20 = -63.208694
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111000000110011111110010001000;
		b = 32'b00101111000010100111110100001010;
		correct = 32'b01100111101001101001101010101111;
		#400 //1.2492865e+34 * 1.259545e-10 = 1.5735325e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100011101111111110010000110000;
		b = 32'b11100110001011011101111001111010;
		correct = 32'b11001010100000100101001111111000;
		#400 //2.0804903e-17 * -2.0526834e+23 = -4270588.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110101011011000010010110010;
		b = 32'b11100100110000000010000000101100;
		correct = 32'b11100100000000100011100101010100;
		#400 //0.338903 * -2.8352745e+22 = -9.608831e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101001001111110111001000101011;
		b = 32'b00001000101010011000111111110101;
		correct = 32'b00110010011111011001110000001101;
		#400 //1.4465248e+25 * 1.0205162e-33 = 1.476202e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111011001100000101001000100000;
		b = 32'b10101101111100001000111100101101;
		correct = 32'b00101001101001011010111110011011;
		#400 //-0.002690442 * -2.7348424e-11 = 7.3579347e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010010000000101011000101111101;
		b = 32'b11010101011100111000000010000100;
		correct = 32'b10100111111110001010000000101100;
		#400 //4.123954e-28 * -16733331000000.0 = -6.9007486e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011111010011001000010101110;
		b = 32'b10011000110011100100011000010100;
		correct = 32'b00100101001111000011001001011100;
		#400 //-30613852.0 * -5.3320513e-24 = 1.6323463e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001001000111010010100101110100;
		b = 32'b01100101111001111111000101101000;
		correct = 32'b11101111100011100110010010011100;
		#400 //-643735.25 * 1.3691498e+23 = -8.8137e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110101011010110101111110001011;
		b = 32'b00010111110000100101100101100100;
		correct = 32'b10001101101100101011000010010111;
		#400 //-8.7683355e-07 * 1.2559522e-24 = -1.1012609e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011100010101000011101110110011;
		b = 32'b11001111100111000111101001101101;
		correct = 32'b10101100100000011011100111100000;
		#400 //7.0222075e-22 * -5250538000.0 = -3.687037e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001110110101010000101100100001;
		b = 32'b10010000001100110001100010001001;
		correct = 32'b00011111100101010000101100110011;
		#400 //-1787138200.0 * -3.5320427e-29 = 6.312248e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011111110101100011110111000100;
		b = 32'b10101101000011010110101011011000;
		correct = 32'b00001101011011001011001011011111;
		#400 //-9.073471e-20 * -8.038646e-12 = 7.2938423e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001001101101110010100111110011;
		b = 32'b11000001001011011010101011100011;
		correct = 32'b11001011011110001000001100111011;
		#400 //1500478.4 * -10.85422 = -16286523.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001110101100000100000110010010;
		b = 32'b11001100110001000111011110011111;
		correct = 32'b10011100000001110100010010010000;
		#400 //4.345049e-30 * -103005430.0 = -4.475637e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001100101100000000010010001000;
		b = 32'b11100111111001111100001000101110;
		correct = 32'b11110101000111110101100110011010;
		#400 //92283970.0 * -2.1888973e+24 = -2.0200013e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100001110001111011111111101110;
		b = 32'b10111101001000111101111111011101;
		correct = 32'b01011111011111111011101111000010;
		#400 //-4.605915e+20 * -0.040008415 = 1.8427536e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100001001101111010111111111000;
		b = 32'b00110001010011011000010111001110;
		correct = 32'b01010011000100110111011111101100;
		#400 //2.1177713e+20 * 2.9907485e-09 = 633372150000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001100010001101000110110100010;
		b = 32'b01000011111001100101111011001111;
		correct = 32'b10010000101100101010110011001000;
		#400 //-1.5295986e-31 * 460.7407 = -7.047483e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111111011100011110011110101100;
		b = 32'b00001111101101100101110010100010;
		correct = 32'b00001111101011000101001000111101;
		#400 //0.9449413 * 1.7982266e-29 = 1.6992186e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100000101011100101101110110111;
		b = 32'b01000000000001010110010001000011;
		correct = 32'b00100001001101011011001111011111;
		#400 //2.9537438e-19 * 2.0842445 = 6.1563243e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011100100011110110010001011101;
		b = 32'b01111000111101001100001111100110;
		correct = 32'b01010110000010010001100101100011;
		#400 //9.48889e-22 * 3.971543e+34 = 37685530000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000011101011100110111100011010;
		b = 32'b01000011110101101011001000000011;
		correct = 32'b00001000000100100100101000101011;
		#400 //1.02523085e-36 * 429.39072 = 4.402246e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000001100100011100011101000011;
		b = 32'b01010000010110010101101011000110;
		correct = 32'b01010010011101111000101100110001;
		#400 //18.222296 * 14586419000.0 = 265798040000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100011101110101111101110010101;
		b = 32'b10011100110110000111100110111101;
		correct = 32'b01000001000111100001110100110001;
		#400 //-6.8984456e+21 * -1.432515e-21 = 9.882127
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011010010110110111110001101000;
		b = 32'b11011101001101000011101011100101;
		correct = 32'b00111000000110101000010111111000;
		#400 //-4.5388633e-23 * -8.11684e+17 = 3.684123e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111000111100001010111011000011;
		b = 32'b00101111001001101011100010100111;
		correct = 32'b10101000100111001011111011101101;
		#400 //-0.00011476644 * 1.5163214e-10 = -1.740228e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110011101000011101000011011100;
		b = 32'b10111100111110011100101001000000;
		correct = 32'b01110001000111011110001111111101;
		#400 //-2.5640746e+31 * -0.030491948 = 7.818363e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011001010000100101011000110001;
		b = 32'b00110111111111110110111001001101;
		correct = 32'b01010001110000011110011110010110;
		#400 //3418807000000000.0 * 3.0449732e-05 = 104101760000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110111100111001111011010001;
		b = 32'b10001011000010110010111011011001;
		correct = 32'b00000010100001000111001111010001;
		#400 //-7.260453e-06 * -2.680567e-32 = 1.9462132e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111100000101011001110001011011;
		b = 32'b10001010010100000100110100001000;
		correct = 32'b00000110111100110111100000011101;
		#400 //-0.009131516 * -1.0029324e-32 = 9.158293e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101000011000000100010101001000;
		b = 32'b00100010101000010111100110000110;
		correct = 32'b10001011100011010111011000001000;
		#400 //-1.2449521e-14 * 4.3767805e-18 = -5.448882e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001010101000011111100111100100;
		b = 32'b00001001011010011110111100011011;
		correct = 32'b10010100100101000000001110111010;
		#400 //-5307634.0 * 2.8158782e-33 = -1.4945651e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110110001101111110000000100111;
		b = 32'b11101000100011100111101110011101;
		correct = 32'b11011111010011001010111000111110;
		#400 //2.7399599e-06 * -5.3828504e+24 = -1.4748794e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111110010010000100000111100001;
		b = 32'b10001000111110001011110111001110;
		correct = 32'b01000111110000101001010001001100;
		#400 //-6.6546915e+37 * -1.497058e-33 = 99624.59
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101011100011101100010011000100;
		b = 32'b00100101011011111000011110011001;
		correct = 32'b10010001100001011001010101010010;
		#400 //-1.014432e-12 * 2.0775888e-16 = -2.1075726e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010111010011010111111001101001;
		b = 32'b11000001010010100100100001100011;
		correct = 32'b11011001001000100101111111011010;
		#400 //225942810000000.0 * -12.642673 = -2856521000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101101011101010100100010110001;
		b = 32'b10011110010000000110100110001100;
		correct = 32'b11001100001110000101101110100110;
		#400 //4.7444816e+27 * -1.0186222e-20 = -48328344.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000110110110010000010110111100;
		b = 32'b01011101000100110010101000101000;
		correct = 32'b01100100011110011000010000010000;
		#400 //27778.867 * 6.627708e+17 = 1.8411022e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000001110000001000010010000101;
		b = 32'b01001011001100101000100111111111;
		correct = 32'b11001101100001100100001111101011;
		#400 //-24.064707 * 11700735.0 = -281574750.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110110010010110001101011110011;
		b = 32'b10011000100010001010001010110001;
		correct = 32'b11001111010110001100111011001001;
		#400 //1.0298661e+33 * -3.5319452e-24 = -3637430500.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001101100101111100111011101110;
		b = 32'b01100001000110110110000111000000;
		correct = 32'b01101111001110000100100010000011;
		#400 //318365120.0 * 1.7914306e+20 = 5.7032903e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100011011110001000101111101001;
		b = 32'b00101011000011010010110111011101;
		correct = 32'b00001111000010010001000110010110;
		#400 //1.3473734e-17 * 5.015691e-13 = 6.7580084e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000010110011011011001001100001;
		b = 32'b01101001100011010110111111100100;
		correct = 32'b10101100111000110100101001001110;
		#400 //-3.0224427e-37 * 2.1373366e+25 = -6.4599775e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010000001000010100011101001;
		b = 32'b11010100101100010111111001010001;
		correct = 32'b01001111001101110100001011111110;
		#400 //-0.00050414965 * -6098627600000.0 = 3074621000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101010011000001110111100000111;
		b = 32'b00100010111000001101101101001010;
		correct = 32'b11001101110001011001000111010100;
		#400 //-6.798204e+25 * 6.0947503e-18 = -414333570.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110001110011110010111010110000;
		b = 32'b10011111010101000110100100001100;
		correct = 32'b11010001101010111110011110101110;
		#400 //2.0518348e+30 * -4.497964e-20 = -92290790000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111000110011101010101001110110;
		b = 32'b00101000111010011000001001000011;
		correct = 32'b10100010001111001000001001001110;
		#400 //-9.854596e-05 * 2.5924688e-14 = -2.5547734e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101111010000100001111000111110;
		b = 32'b00101101100101011111011001101010;
		correct = 32'b11011101011000110110110011100111;
		#400 //-6.0076652e+28 * 1.7048769e-11 = -1.02423295e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100011111010100100110001001010;
		b = 32'b10111110111111010100000011110000;
		correct = 32'b11100011011001111100100011010100;
		#400 //8.6440706e+21 * -0.49463606 = -4.275669e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011110001100100011111011101011;
		b = 32'b01001100101001000010111110001010;
		correct = 32'b01101011011001001010001011010000;
		#400 //3.2109904e+18 * 86080590.0 = 2.7640395e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100111000101000000010111100111;
		b = 32'b10111010000000011101101111101010;
		correct = 32'b00100001100101100010110001000100;
		#400 //-2.0542326e-15 * -0.0004953729 = 1.0176112e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011010000100001101101101100000;
		b = 32'b00111110101000001111010100111010;
		correct = 32'b11011001001101100010011110111110;
		#400 //-1.01934e+16 * 0.31437093 = -3204509000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100110111000101000100110000000;
		b = 32'b00100100001100100001011111101100;
		correct = 32'b10001011100111011001100011000110;
		#400 //-1.571917e-15 * 3.861786e-17 = -6.070407e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101110111110010111011101011101;
		b = 32'b00110001011011111101010101011011;
		correct = 32'b11100000111010011011011001011001;
		#400 //-3.8603034e+28 * 3.4900356e-09 = -1.3472597e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111001000001010110101010001010;
		b = 32'b11000000111010010000011001010101;
		correct = 32'b11111010011100101110001010001001;
		#400 //4.329602e+34 * -7.282023 = -3.1528263e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110001110111000010100110100011;
		b = 32'b10100001111100000001011001110011;
		correct = 32'b11010100010011100111101001010111;
		#400 //2.1803852e+30 * -1.6268975e-18 = -3547263100000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011001110111100010110011111010;
		b = 32'b00011010110010100000111010000010;
		correct = 32'b10110101001011110101110000010101;
		#400 //-7817112000000000.0 * 8.356868e-23 = -6.532658e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111100000110101110111101011011;
		b = 32'b00110100001000111000000011101001;
		correct = 32'b11110000110001011110100011010111;
		#400 //-3.2178737e+36 * 1.5227455e-07 = -4.9000026e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111110001100000010111010100000;
		b = 32'b10101010111100110010010001010110;
		correct = 32'b11101001101001110101010101000100;
		#400 //5.8546555e+37 * -4.3190684e-13 = -2.5286658e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000101010101100000100001100110;
		b = 32'b11100011101101000001100011110010;
		correct = 32'b11101001100101101001001011000011;
		#400 //3424.525 * -6.644423e+21 = -2.2753992e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010001000001110101110000010000;
		b = 32'b11000101010010011001010111010011;
		correct = 32'b00010110110101010010110100000001;
		#400 //-1.0677991e-28 * -3225.364 = 3.4440407e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111000111111001001011000001100;
		b = 32'b10010100100011111011010001101101;
		correct = 32'b10001110000011011100100111010110;
		#400 //0.00012044245 * -1.4510475e-26 = -1.7476772e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010001011111000111010011001110;
		b = 32'b00110011101011101011100110100111;
		correct = 32'b00000101101011000100111001111001;
		#400 //1.9915288e-28 * 8.1362764e-08 = 1.6203629e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001100011010001101111100000010;
		b = 32'b01110000011001101110001010011011;
		correct = 32'b11111101010100100000011001111110;
		#400 //-61045770.0 * 2.85822e+29 = -1.7448224e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001011000101000000110001001001;
		b = 32'b00111011010101011110010011000011;
		correct = 32'b10000110111101110110010100001001;
		#400 //-2.8513006e-32 * 0.0032637573 = -9.305953e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110001001010001111011010000111;
		b = 32'b00000101101000100000011011010000;
		correct = 32'b10110111010101011110000100000001;
		#400 //-8.3666424e+29 * 1.523691e-35 = -1.2748177e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110010101101011101110010010110;
		b = 32'b00010000110011011111001000100010;
		correct = 32'b11000100000100100100110110100111;
		#400 //-7.204283e+30 * 8.123131e-29 = -585.2133
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000001101110010010010001000101;
		b = 32'b10010111000010111011100011111011;
		correct = 32'b00011001010010100001100011110010;
		#400 //-23.14271 * -4.51468e-25 = 1.0448193e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000000110001000010011101010000;
		b = 32'b01001000110101001101001001010100;
		correct = 32'b10001010001000110001000110110111;
		#400 //-1.801386e-38 * 435858.62 = -7.851496e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011101101100010010000101010000;
		b = 32'b10100000111010101111101111000000;
		correct = 32'b00111111001000101001011010100100;
		#400 //-1.5954463e+18 * -3.9807736e-19 = 0.6351111
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001101110001110011010100100011;
		b = 32'b11010101000001101001101100011000;
		correct = 32'b11100011010100010111110100000000;
		#400 //417768540.0 * -9250043000000.0 = -3.8643767e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110101110000001010100000101;
		b = 32'b01111100010010001010110000011100;
		correct = 32'b01111011100100000100110000101110;
		#400 //0.35953537 * 4.1678007e+36 = 1.4984717e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111001111101000011100100100001;
		b = 32'b11101011011101110111110001110110;
		correct = 32'b11100101111011000001100111011011;
		#400 //0.0004658187 * -2.9919243e+26 = -1.3936943e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000001001111001000110011000011;
		b = 32'b10000100011001011101011000101101;
		correct = 32'b00000110001010010100011110101001;
		#400 //-11.784366 * -2.7017165e-36 = 3.1838015e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000010101101100101010001111010;
		b = 32'b10001101000001000110100100010101;
		correct = 32'b10010000001111001001110011001101;
		#400 //91.16499 * -4.080213e-31 = -3.7197257e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111000000001011111010110100010;
		b = 32'b01111011111000110100100111001110;
		correct = 32'b01110100011011011101111011011011;
		#400 //3.1938434e-05 * 2.3602966e+36 = 7.538418e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000001011110111110110001001111;
		b = 32'b11000010101110011001011001001111;
		correct = 32'b01000100101101101010000110101111;
		#400 //-15.745193 * -92.79357 = 1461.0526
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000110010000101100010010100010;
		b = 32'b10001111010010101111100111100010;
		correct = 32'b10010110000110100110110101000101;
		#400 //12465.158 * -1.00074946e-29 = -1.24745e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110000011111110010011110101000;
		b = 32'b10110001000000101000000101011111;
		correct = 32'b10100010000000100001001100010101;
		#400 //9.2824815e-10 * -1.8991029e-09 = -1.7628387e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001000100000111111001110100001;
		b = 32'b01001111110011011111110110000110;
		correct = 32'b00011000110101000101100110001010;
		#400 //7.941553e-34 * 6911888400.0 = 5.4891127e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010101110111011100011011101001;
		b = 32'b01000011100100110000001110111010;
		correct = 32'b10011001111111101011100011100101;
		#400 //-8.9575014e-26 * 294.0291 = -2.6337663e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011101001001101011100000011010;
		b = 32'b10010110011001111100111001001000;
		correct = 32'b00110100000101101111011001110110;
		#400 //-7.508363e+17 * -1.8725122e-25 = 1.40595e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100100111001010100101000100010;
		b = 32'b11111001111001111010110000101111;
		correct = 32'b11011111010011111000000000011101;
		#400 //9.9438505e-17 * -1.5036411e+35 = -1.4951983e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010001001110101011001011100010;
		b = 32'b10001010110111000101011000010111;
		correct = 32'b10011100101000001011000010000011;
		#400 //50116567000.0 * -2.1217613e-32 = -1.0633539e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010011101110000000001100111011;
		b = 32'b11101000111001001101101101101111;
		correct = 32'b01111101001001001000000010011011;
		#400 //-1580656400000.0 * -8.645979e+24 = 1.3666322e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001000111100110001111100011011;
		b = 32'b01001001111100111101110111011001;
		correct = 32'b10010011011001111001100100110111;
		#400 //-1.4632343e-33 * 1997755.1 = -2.923184e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110101010010001011001011111010;
		b = 32'b01100010100110110111011011100011;
		correct = 32'b11011000011100111100001100100100;
		#400 //-7.476625e-07 * 1.433906e+21 = -1072077800000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110011001010001011100011111000;
		b = 32'b01010001110110100011001011110101;
		correct = 32'b11000101100011111100111100011001;
		#400 //-3.9283776e-08 * 117144720000.0 = -4601.887
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010000101000001111100111001101;
		b = 32'b01010010111101001100001111111001;
		correct = 32'b10100100000110011110100101010010;
		#400 //-6.349375e-29 * 525629950000.0 = -3.3374216e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100000100011111010001000000011;
		b = 32'b00001111010001110111001001110111;
		correct = 32'b10110000010111111100111001010010;
		#400 //-8.2798706e+19 * 9.833503e-30 = -8.1420126e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100010110111001010011000111101;
		b = 32'b01001001101001101010101001010001;
		correct = 32'b00101101000011111010011010011000;
		#400 //5.980713e-18 * 1365322.1 = 8.1656e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001101001000101000110101110101;
		b = 32'b11101011100001111100101001000001;
		correct = 32'b00111001001011000111001000001011;
		#400 //-5.0090377e-31 * -3.283202e+26 = 0.00016445683
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100101011111111111000100000110;
		b = 32'b01000110100000001011110100101001;
		correct = 32'b00101100100000001011010110100001;
		#400 //2.2199386e-16 * 16478.58 = 3.6581437e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101111000110110101100011111101;
		b = 32'b01100010110010011111100001000101;
		correct = 32'b01010010011101010001111100001101;
		#400 //1.4128783e-10 * 1.8628426e+21 = 263196980000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111101011010111001101010111000;
		b = 32'b11100000000110010000011101010110;
		correct = 32'b11011110000011001101011000111000;
		#400 //0.0575206 * -4.4107507e+19 = -2.53709e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010001110101111111011000100110;
		b = 32'b11010010010111101110100101110000;
		correct = 32'b10100100101111000000110001100010;
		#400 //3.407272e-28 * -239349800000.0 = -8.155298e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000011101101001010000010101010;
		b = 32'b11111000101101001000001111001010;
		correct = 32'b11111100111111101011101111101001;
		#400 //361.2552 * -2.92902e+34 = -1.05812374e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011101110100100101011111010110;
		b = 32'b11010011000001111111011010111001;
		correct = 32'b01110001010111110110111000010101;
		#400 //-1.8946023e+18 * -583959900000.0 = 1.1063718e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010000111101001110101001011110;
		b = 32'b10101011110100000111001011000000;
		correct = 32'b10111101010001110110110000110100;
		#400 //32872002000.0 * -1.4811138e-12 = -0.048687175
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101101000100100001001011001000;
		b = 32'b01001011100101101100000010011111;
		correct = 32'b10111001001011000000100111010100;
		#400 //-8.303309e-12 * 19759422.0 = -0.0001640686
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101101000101100110100010010101;
		b = 32'b10100010111010100011011111100011;
		correct = 32'b00010000100010011001110001101110;
		#400 //-8.549735e-12 * -6.3485e-18 = 5.427799e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001000000111100001101000001100;
		b = 32'b01101100011000010011011111000110;
		correct = 32'b01110101000010110001011101010110;
		#400 //161896.19 * 1.0890868e+27 = 1.7631899e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011000011110110001001100100100;
		b = 32'b11110001111000100111010111000101;
		correct = 32'b11001010110111100001101001100111;
		#400 //3.2450653e-24 * -2.2427516e+30 = -7277875.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000111000110011111110001110101;
		b = 32'b11100101001011101111011110011010;
		correct = 32'b10101100110100100111110100001101;
		#400 //1.1584631e-34 * -5.16412e+22 = -5.9824424e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010011101011010001010011010001;
		b = 32'b00001101100001101100000010001101;
		correct = 32'b10100001101101100011011000101001;
		#400 //-1486757200000.0 * 8.3047425e-31 = -1.2347136e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000000010000011010001101011000;
		b = 32'b01100101101001010100111010100000;
		correct = 32'b00100110001010011000100111000010;
		#400 //6.027904e-39 * 9.758011e+22 = 5.882035e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110110010011011010000111000110;
		b = 32'b00000010000011100000111001000100;
		correct = 32'b00111000111001000011011001100011;
		#400 //1.04267775e+33 * 1.0436606e-37 = 0.000108820175
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010000011100100000111111011111;
		b = 32'b01110001110011101111101110010011;
		correct = 32'b01000010110000111011011010100110;
		#400 //4.773831e-29 * 2.0498575e+30 = 97.856735
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110100101101110110101001111000;
		b = 32'b00010000100001010110000011010101;
		correct = 32'b01000101101111110001111101100010;
		#400 //1.1625363e+32 * 5.2608444e-29 = 6115.923
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101010010010000101110000110101;
		b = 32'b00011100100100111110001001011011;
		correct = 32'b10000111011001110111110000110110;
		#400 //-1.7795559e-13 * 9.786156e-22 = -1.7415011e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110011010100000000011011001;
		b = 32'b00101110100111011100001010001111;
		correct = 32'b00101101100100000011010001011100;
		#400 //0.22851886 * 7.174094e-11 = 1.6394157e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111010000111110100001011111110;
		b = 32'b10011101000100011000110000100000;
		correct = 32'b01010111101101010001100000111101;
		#400 //-2.067335e+35 * -1.9263033e-21 = 398231400000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110101110100111110010010001010;
		b = 32'b11001110111101010100010010110100;
		correct = 32'b01000101010010110000001010010110;
		#400 //-1.5787239e-06 * -2057460200.0 = 3248.1616
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011001110101100010011110111110;
		b = 32'b11110111100100000010000000100110;
		correct = 32'b01010001111100010010001001111111;
		#400 //-2.2143133e-23 * -5.846428e+33 = 129458230000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111001100100100001011000100100;
		b = 32'b11000011111100111011011110111101;
		correct = 32'b00111110000010110001001111011110;
		#400 //-0.00027863786 * -487.43546 = 0.13581797
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011110110110111010000010100011;
		b = 32'b10111110001000001001001000100101;
		correct = 32'b11011101100010011100000111000111;
		#400 //7.912914e+18 * -0.1568075 = -1.2408042e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010000100101000101100010000010;
		b = 32'b10011110100001010000000111111110;
		correct = 32'b10101111100110100010011001000110;
		#400 //19910627000.0 * -1.4082747e-20 = -2.8039632e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100000011111011101110000101010;
		b = 32'b11100111100011111011100110101100;
		correct = 32'b01001000100011101000011000011010;
		#400 //-2.150278e-19 * -1.3574469e+24 = 291888.8
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101000000001101100100011011100;
		b = 32'b00110101010011000010110101010110;
		correct = 32'b00011101110101101111111111011100;
		#400 //7.482049e-15 * 7.6061895e-07 = 5.690988e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001010100011100010111001110000;
		b = 32'b00011001110101110010110100111001;
		correct = 32'b10100100111011110000010000111100;
		#400 //-4659000.0 * 2.2248744e-23 = -1.036569e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111100001100101111001011000111;
		b = 32'b00110000010001100000000111000101;
		correct = 32'b11101101000010100110100100000011;
		#400 //-3.7166118e+36 * 7.2034495e-10 = -2.6772427e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011101000010101100011100101110;
		b = 32'b10111101011100111101000000010110;
		correct = 32'b11011011000001000010101111011110;
		#400 //6.2500075e+17 * -0.059524618 = -3.720293e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010000001110000100000010000101;
		b = 32'b11001000011101011101100001100100;
		correct = 32'b00011001001100001111000101111110;
		#400 //-3.6337306e-29 * -251745.56 = 9.147756e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010111101101110110011001111010;
		b = 32'b01110100001011000000010001010110;
		correct = 32'b01001100011101100111011111101010;
		#400 //1.1851967e-24 * 5.4514343e+31 = 64610216.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001011000101001111100000000011;
		b = 32'b10010010100100000000110100010100;
		correct = 32'b10011110001001111010011000111100;
		#400 //9762819.0 * -9.090902e-28 = -8.875283e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110111110101000101010111110;
		b = 32'b00101110110111111000011110000010;
		correct = 32'b10100110010110101100001101111010;
		#400 //-7.4667323e-06 * 1.0164937e-10 = -7.5898864e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010110011111110001110111101000;
		b = 32'b00110101100100110111111110111011;
		correct = 32'b01001100100100101111110101110110;
		#400 //70125978000000.0 * 1.0989528e-06 = 77065140.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001111000001110101100000000110;
		b = 32'b11010000110101011010010110011111;
		correct = 32'b01100000011000011110011110011010;
		#400 //-2270692900.0 * -28675210000.0 = 6.5112595e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001100100111010001001111000011;
		b = 32'b00100000110000101000000010010010;
		correct = 32'b00101101111011101010111110111010;
		#400 //82353690.0 * 3.294996e-19 = 2.7135506e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100011000001101111100100110101;
		b = 32'b11100001110010011010000001111000;
		correct = 32'b11000101010101001001110010001011;
		#400 //7.316926e-18 * -4.6491982e+20 = -3401.784
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111110001111010100010011011000;
		b = 32'b00001011001011001110110000111101;
		correct = 32'b01001001111111111011000111010011;
		#400 //6.2895387e+37 * 3.330372e-32 = 2094650.4
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011000000101100101010101010001;
		b = 32'b10101100001010110011010110110110;
		correct = 32'b01000100110010010001010100001111;
		#400 //-661172700000000.0 * -2.4330377e-12 = 1608.6581
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100001100010000000010001000111;
		b = 32'b10001000101011001101010001011010;
		correct = 32'b00101010101101111010011101100110;
		#400 //-3.1363318e+20 * -1.0401797e-33 = 3.2623486e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000010010111100110001011000;
		b = 32'b01001010110110111101001000011000;
		correct = 32'b10111011101011101111111100010000;
		#400 //-7.414136e-10 * 7203084.0 = -0.0053404644
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011100110101111001101101010010;
		b = 32'b10100100110111110001011100101010;
		correct = 32'b11000010001110111110001111001111;
		#400 //4.8550317e+17 * -9.6750075e-17 = -46.97247
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010100110001010011110100000;
		b = 32'b11010011010010001100111110101011;
		correct = 32'b01001110011011110111110110010101;
		#400 //-0.0011646636 * -862477550000.0 = 1004496200.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110000110111110010010011111101;
		b = 32'b01101110100111001110110101100010;
		correct = 32'b01100000000010001100100101110101;
		#400 //1.6235898e-09 * 2.428332e+28 = 3.942615e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010000100000110001000011100110;
		b = 32'b10001101110110001000000010101000;
		correct = 32'b10011110110111011011000001000001;
		#400 //17591382000.0 * -1.3343001e-30 = -2.3472182e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000111000011000011001110111110;
		b = 32'b01000101011100000000011101110111;
		correct = 32'b10001101000000110111010010011001;
		#400 //-1.0547635e-34 * 3840.4666 = -4.050784e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100100000010000110010010100011;
		b = 32'b11110100110000100110000100100111;
		correct = 32'b11011001010011110010000000001101;
		#400 //2.9575542e-17 * -1.2320265e+32 = -3643785000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000010001101100001100000011101;
		b = 32'b11011010100001100010010110101110;
		correct = 32'b00011101001111101101011011011001;
		#400 //-1.3378168e-37 * -1.8879538e+16 = 2.5257364e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010011101101010010100010001011;
		b = 32'b10111110111010111110101011100111;
		correct = 32'b01010011001001101111001001110010;
		#400 //-1556138600000.0 * -0.46077654 = 717032100000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111110010110111001101110100100;
		b = 32'b11011100011110101000000110101101;
		correct = 32'b01011011010101101110010100111100;
		#400 //-0.21446091 * -2.820453e+17 = 6.048769e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101000110010010101100010001111;
		b = 32'b00110111110111001111001000100100;
		correct = 32'b11100001001011011100011010001101;
		#400 //-7.606634e+24 * 2.63388e-05 = -2.0034961e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010010000010110011000100111001;
		b = 32'b10011100011111010000111001000111;
		correct = 32'b00101111000010011001011101101001;
		#400 //-149456570000.0 * -8.372913e-22 = 1.2513869e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100010111111100000000000001111;
		b = 32'b10011111111110111101101001010101;
		correct = 32'b10000011011110011110001010101111;
		#400 //6.88469e-18 * -1.06663835e-19 = -7.3434743e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101000111000011101010010110100;
		b = 32'b01001101101011011101111101011010;
		correct = 32'b00110111000110010110000111000101;
		#400 //2.5072263e-14 * 364637000.0 = 9.142274e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101100010101110111000111000111;
		b = 32'b01110100111110110001110111000101;
		correct = 32'b11100001110100110101010110011100;
		#400 //-3.0616497e-12 * 1.5916386e+32 = -4.8730398e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110101011001101101100101010011;
		b = 32'b01011010111111011010110110100011;
		correct = 32'b11010000111001001100000101011011;
		#400 //-8.5997925e-07 * 3.5702042e+16 = -30703016000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001101100100110011110101100000;
		b = 32'b00110001101111100011011000010101;
		correct = 32'b10111111110110101100110101010001;
		#400 //-308784130.0 * 5.535876e-09 = -1.7093908
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010110101001100000100010010110;
		b = 32'b10010100100010001111111010001111;
		correct = 32'b00101011101100011011001101010010;
		#400 //-91277900000000.0 * -1.3832896e-26 = 1.2626378e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111111000001110010101000010;
		b = 32'b11000001010101001100001010000100;
		correct = 32'b11001001101110101110100010111100;
		#400 //115146.516 * -13.297489 = -1531159.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001111010011100000011011101100;
		b = 32'b01000111010001000111010100001001;
		correct = 32'b10010111000111100001101101111101;
		#400 //-1.0157917e-29 * 50293.035 = -5.108725e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011111101000011110111011100101;
		b = 32'b00010001110100000000101000000111;
		correct = 32'b00110010000000111001100001110010;
		#400 //2.333703e+19 * 3.2822793e-28 = 7.659866e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110100111111000011101101001;
		b = 32'b10100111100101111110011011001011;
		correct = 32'b10100110101111010101000101100010;
		#400 //0.31157997 * -4.2161145e-15 = -1.3136568e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110101000110101000111000010110;
		b = 32'b01110001111101001010110110110011;
		correct = 32'b01100111100100111011100001001011;
		#400 //5.7576233e-07 * 2.4231786e+30 = 1.395175e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111010001110101010100001100000;
		b = 32'b00100100111011110000011011101001;
		correct = 32'b11011111101011100100100000111011;
		#400 //-2.4229557e+35 * 1.03661434e-16 = -2.5116705e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111001010011100111011100011111;
		b = 32'b01101100101101101101101101010110;
		correct = 32'b11100110100100110111100110010101;
		#400 //-0.00019690067 * 1.7684823e+27 = -3.4821533e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111110011100110100111110111110;
		b = 32'b00001111011010110100100001101100;
		correct = 32'b10001110010111111001111100001000;
		#400 //-0.23760888 * 1.16003425e-29 = -2.7563443e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010001111100100011100110011011;
		b = 32'b01111101101110011101010101110001;
		correct = 32'b01010000001011111101010110010110;
		#400 //3.821637e-28 * 3.087693e+37 = 11800041000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110011111111011101100000100;
		b = 32'b10100111110000001100101011111111;
		correct = 32'b00011110110000001001011100001011;
		#400 //-3.8106818e-06 * -5.3510794e-15 = 2.039126e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010111001011010110011101001001;
		b = 32'b01111111111101100110000010000010;
		correct = 32'b01111111111101100110000010000010;
		#400 //190659120000000.0 * nan = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000000100011011001100101110011;
		b = 32'b01110110010100010010111000001100;
		correct = 32'b11110111011001110110011101111110;
		#400 //-4.4249816 * 1.06066795e+33 = -4.693436e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111100111000101100111100011001;
		b = 32'b10101111110011101110011100101001;
		correct = 32'b10101101001101110100111101110011;
		#400 //0.027686642 * -3.763543e-10 = -1.0419987e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001011010000100001000110010110;
		b = 32'b11000110010110110010100111111101;
		correct = 32'b00010010001001100010010011100000;
		#400 //-3.737627e-32 * -14026.497 = 5.2425816e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010001011100011011000110111111;
		b = 32'b10011111010101011111111100100111;
		correct = 32'b00110001010010100000100111001001;
		#400 //-64879325000.0 * -4.531556e-20 = 2.940043e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100101000111010111111010101001;
		b = 32'b11001000100110110000110100110000;
		correct = 32'b11101110001111101100011110011011;
		#400 //4.648425e+22 * -317545.5 = -1.4760865e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101000000000010111101010000001;
		b = 32'b10110110000100011000110010001011;
		correct = 32'b11011110100100110011101011110001;
		#400 //2.4457803e+24 * -2.168849e-06 = -5.3045284e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111101010101101010111110110100;
		b = 32'b00100111000100101011011111011010;
		correct = 32'b11100100111101100001010011000110;
		#400 //-1.7835443e+37 * 2.0361236e-15 = -3.6315167e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010100100101100001110110110010;
		b = 32'b10000001011010001100010000000011;
		correct = 32'b00010110100010000111110111011010;
		#400 //-5157946400000.0 * -4.2752302e-38 = 2.2051409e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101101010011011010011001000010;
		b = 32'b10100100001101110100011110100101;
		correct = 32'b01010010000100110011101101100111;
		#400 //-3.9778388e+27 * -3.9742485e-17 = 158089200000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100001000001111101001000110011;
		b = 32'b00100110011011000011100010100100;
		correct = 32'b10000111111110101010011110101000;
		#400 //-4.6017976e-19 * 8.195571e-16 = -3.7714359e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010001111110011011001110110001;
		b = 32'b11011111001101110111001001010101;
		correct = 32'b11110001101100101110111011111000;
		#400 //134057700000.0 * -1.3218721e+19 = -1.7720713e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110110010001011101111111011100;
		b = 32'b10011110101110100010000010111011;
		correct = 32'b10010101100011111101110111110010;
		#400 //2.948559e-06 * -1.9707053e-20 = -5.810741e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100011100100011111011111110100;
		b = 32'b11000111111101001111010001101011;
		correct = 32'b10101100000010111010101110110010;
		#400 //1.5825944e-17 * -125416.836 = -1.9848398e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010101100111110011010101100100;
		b = 32'b01100111111011111100100000001100;
		correct = 32'b11111110000101010001111101000010;
		#400 //-21881457000000.0 * 2.2646716e+24 = -4.955432e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110101010011101010001111011100;
		b = 32'b01111101110111110100101011000100;
		correct = 32'b01110011101101000011110100010110;
		#400 //7.6979427e-07 * 3.7100756e+37 = 2.855995e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101000001000100110000101110101;
		b = 32'b11001001000000010010101100100101;
		correct = 32'b00110001101000111101110011110100;
		#400 //-9.013939e-15 * -529074.3 = 4.769044e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111111000000100110011011100101;
		b = 32'b00101001001100010011110000000001;
		correct = 32'b00101000101101001000111101101010;
		#400 //0.50938255 * 3.935394e-14 = 2.004621e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001010100111001010110011101110;
		b = 32'b10111000110000000011011100110001;
		correct = 32'b10000011111010110100011011110011;
		#400 //1.5087302e-32 * -9.165554e-05 = -1.3828348e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010100001101001010100011001011;
		b = 32'b10111100111010011011111001010010;
		correct = 32'b01010001101001001111001111110000;
		#400 //-3103704000000.0 * -0.028533135 = 88558400000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001101011110100001001101101010;
		b = 32'b10110100111010001111011000100111;
		correct = 32'b10000010111000111001001000001101;
		#400 //7.7060567e-31 * -4.3392467e-07 = -3.3438481e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010101010110000111100111010;
		b = 32'b01001111010010001001100101110000;
		correct = 32'b11001010100001100000101001101100;
		#400 //-0.0013050803 * 3365499000.0 = -4392246.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111001011101001010110110110110;
		b = 32'b00111101011000100010001110110000;
		correct = 32'b11110111010110000010001101110111;
		#400 //-7.940273e+34 * 0.055209816 = -4.3838103e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110010011110101100000001101001;
		b = 32'b10111010010111011110001100010110;
		correct = 32'b10101101010110010101011010001001;
		#400 //1.4595664e-08 * -0.00084643194 = -1.23542366e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000010000110010010010101011001;
		b = 32'b11001000011000100011100000010101;
		correct = 32'b00001011000001110101010010000101;
		#400 //-1.1251383e-37 * -231648.33 = 2.606364e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101100011100110001110000000110;
		b = 32'b00010110011011000100011100111001;
		correct = 32'b01000011011000000110000101111000;
		#400 //1.17560524e+27 * 1.9086402e-25 = 224.38074
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010001001011101111011101111100;
		b = 32'b10011010100010001011110111110110;
		correct = 32'b00101100001110101110101010011101;
		#400 //-46967276000.0 * -5.655518e-23 = 2.6562426e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000100100000011000110110001111;
		b = 32'b11110010101100101010000111001111;
		correct = 32'b01110111101101001100110010100000;
		#400 //-1036.4237 * -7.076345e+30 = 7.3340916e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100010001111100000001010111001;
		b = 32'b11000100101111110001110000011010;
		correct = 32'b00100111100011011101100011100100;
		#400 //-2.5751243e-18 * -1528.8782 = 3.9370515e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110111000000011011110011101100;
		b = 32'b00110001101001100111101011011011;
		correct = 32'b00101001001010001011110110001000;
		#400 //7.732986e-06 * 4.845203e-09 = 3.7467886e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100001111011100010001010100001;
		b = 32'b01100111011100010000000000011110;
		correct = 32'b01001001111000000010111010110101;
		#400 //1.6136674e-18 * 1.1380925e+24 = 1836502.6
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100101101000100000100100000011;
		b = 32'b10010101100100101001111100101101;
		correct = 32'b00111011101110011001101111001000;
		#400 //-9.56487e+22 * -5.9220065e-26 = 0.0056643225
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101000111111100101001110111110;
		b = 32'b11100001101101011101011101010101;
		correct = 32'b11001011001101001010011100100010;
		#400 //2.8235982e-14 * -4.1929712e+20 = -11839266.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010111010100100110011110000100;
		b = 32'b10011000111110000000000010001010;
		correct = 32'b10110000110010111101010010111001;
		#400 //231342040000000.0 * -6.410704e-24 = -1.4830653e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001110011000000101010110111100;
		b = 32'b01011110100100000101000000001010;
		correct = 32'b10101101011111001110110010111011;
		#400 //-2.7651411e-30 * 5.199411e+18 = -1.4377106e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000010010011011010100011100001;
		b = 32'b01101101101000100001111011100111;
		correct = 32'b10110000100000100011110110110010;
		#400 //-1.5109487e-37 * 6.271741e+27 = -9.47628e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011010111010110111100101111101;
		b = 32'b00111010001011110101101110100100;
		correct = 32'b01010101101000010100110001010111;
		#400 //3.3140099e+16 * 0.0006689376 = 22168656000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011110100001110000011011011010;
		b = 32'b01110010001100110010111100110100;
		correct = 32'b01010001001111010000010101100000;
		#400 //1.4296515e-20 * 3.5491124e+30 = 50739937000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001111100101101100011100100100;
		b = 32'b01111001101110000000100000001000;
		correct = 32'b01001001110110001100011110111010;
		#400 //1.4867848e-29 * 1.1944319e+35 = 1775863.2
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001110111001010110111100000010;
		b = 32'b01000011111000101010011101011011;
		correct = 32'b11010011010010110010000111111101;
		#400 //-1924628700.0 * 453.30746 = -872448600000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111011001001110001000011001001;
		b = 32'b10001001001010000101101000001101;
		correct = 32'b01000100110110111011101110010001;
		#400 //-8.67454e+35 * -2.0264606e-33 = 1757.8615
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101010000110000011101011001110;
		b = 32'b10100100001000011111000111111011;
		correct = 32'b01001110110000001001100111000000;
		#400 //-4.6008605e+25 * -3.5116275e-17 = 1615650800.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010011111111101000000111100;
		b = 32'b10101111111100110100111101110110;
		correct = 32'b00101010111100110010001000010000;
		#400 //-0.00097585074 * -4.4257903e-10 = 4.3189107e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101000001011101100011110010011;
		b = 32'b10100001110000100111010110101011;
		correct = 32'b10001010100001001100001110010011;
		#400 //9.702216e-15 * -1.3177098e-18 = -1.2784704e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110011111100100110101011000010;
		b = 32'b10110100000011101111101001000110;
		correct = 32'b01101000100001110110010000110110;
		#400 //-3.841251e+31 * -1.331583e-07 = 5.1149443e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011111110011100110010011100001;
		b = 32'b10101111110101011101101100101110;
		correct = 32'b10010000001011000110101010100101;
		#400 //8.7411284e-20 * -3.890021e-10 = -3.4003175e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100100111001100110100100000;
		b = 32'b00100011100010000100011001101111;
		correct = 32'b00101000101001101111000000111010;
		#400 //1254.4102 * 1.477498e-17 = 1.8533884e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101110110001010010111010010011;
		b = 32'b00011110010111111001100010101111;
		correct = 32'b00001101101011000011100100101100;
		#400 //8.966796e-11 * 1.1837096e-20 = 1.0614082e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100100111111010000100111000101;
		b = 32'b01010110111010100100001010001001;
		correct = 32'b11111100011001111000110010110010;
		#400 //-3.7341842e+22 * 128785740000000.0 = -4.809097e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010101001111001011011000001;
		b = 32'b11001010011111000100011101000011;
		correct = 32'b01000101101001010010011100001101;
		#400 //-0.0012786017 * -4133328.8 = 5284.8813
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111110111110100010100000111011;
		b = 32'b11101001001010111000011010010111;
		correct = 32'b01101000101001111001110001100100;
		#400 //-0.48858818 * -1.2960119e+25 = 6.332161e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111011111110100111111101100001;
		b = 32'b00111001010110000101010100111111;
		correct = 32'b01110101110100111010111011100100;
		#400 //2.6013155e+36 * 0.00020631122 = 5.366806e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110100101101001110111011111111;
		b = 32'b10000101000111000100011110111100;
		correct = 32'b10111010010111001110100010101101;
		#400 //1.1468028e+32 * -7.34826e-36 = -0.00084270054
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110000100100100010101111111101;
		b = 32'b11001101101010100000001100000001;
		correct = 32'b10111110110000100010010111011010;
		#400 //1.06354e-09 * -356540450.0 = -0.37919503
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111111110110100010011000011011;
		b = 32'b10010110011001001110100111000011;
		correct = 32'b01111111110110100010011000011011;
		#400 //nan * -1.8491456e-25 = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110110111101000111101000110001;
		b = 32'b10011011000000010101000110000000;
		correct = 32'b01010010011101101111111011001111;
		#400 //-2.4792945e+33 * -1.0696964e-22 = 265209230000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000000110111100010100110000101;
		b = 32'b00000011111111011010010000000011;
		correct = 32'b10000101010111000001110101011110;
		#400 //-6.9425683 * 1.4907659e-36 = -1.0349744e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101111110001101110001011010100;
		b = 32'b10000111010001111100100111001100;
		correct = 32'b00110111100110110011011100011001;
		#400 //-1.231045e+29 * -1.5030399e-34 = 1.8503097e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111110111110011100110100111101;
		b = 32'b00001110000001101000100100100010;
		correct = 32'b10001101100000110100011100111110;
		#400 //-0.48789397 * 1.6582802e-30 = -8.090649e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101110000111111010101110011000;
		b = 32'b10000011110101010011000110101101;
		correct = 32'b10110010100001001111100011000001;
		#400 //1.235389e+28 * -1.253042e-36 = -1.5479943e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000110000011000011011000100001;
		b = 32'b00100000110100110011101111101101;
		correct = 32'b00100111011001110110001011011111;
		#400 //8973.532 * 3.5784446e-19 = 3.2111288e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111010100110001100111000000111;
		b = 32'b00000101001000011010011101101000;
		correct = 32'b11000000010000001111101011111110;
		#400 //-3.9670393e+35 * 7.600931e-36 = -3.0153193
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111010011110011110110001101010;
		b = 32'b10001000101110100110011001110101;
		correct = 32'b10000011101101011111100111001011;
		#400 //0.00095338246 * -1.1218555e-33 = -1.06955735e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001001010001100111110011111000;
		b = 32'b01010010101010100101101110011001;
		correct = 32'b11011100100001000001011000000010;
		#400 //-813007.5 * 365840600000.0 = -2.9743116e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111101000011000111010011001011;
		b = 32'b11010111101010010101011110110001;
		correct = 32'b01010101001110011101001001101110;
		#400 //-0.03429107 * -372388200000000.0 = 12769590000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100000100011001111101011000001;
		b = 32'b11100111000111101101010001000001;
		correct = 32'b11001000001011101110111101001101;
		#400 //2.3882858e-19 * -7.500493e+23 = -179133.2
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100111000101011101000100001101;
		b = 32'b00010101010101101110011001101000;
		correct = 32'b00111100111110111000011100101111;
		#400 //7.074889e+23 * 4.3398714e-26 = 0.030704109
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000000001010010000010110100110;
		b = 32'b10010011011111100101110100010111;
		correct = 32'b10010100001001111111000100010001;
		#400 //2.6409698 * -3.2105204e-27 = -8.478887e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011011000111011100010110110000;
		b = 32'b10101111100110001010011011000011;
		correct = 32'b11001011001111000010100001001110;
		#400 //4.440893e+16 * -2.776713e-10 = -12331086.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111010111011011010011010010101;
		b = 32'b01000100001001101101001000000100;
		correct = 32'b00111111100110101101110011111011;
		#400 //0.001813131 * 667.2815 = 1.2098688
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001101110100100110110101101001;
		b = 32'b01110010001011111111011001110101;
		correct = 32'b11000000100100001010001101100000;
		#400 //-1.2968589e-30 * 3.4853008e+30 = -4.519943
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110110111101011000110101010001;
		b = 32'b00011010110011111110001001000110;
		correct = 32'b00010010010001110110011001001110;
		#400 //7.3180204e-06 * 8.597876e-23 = 6.291943e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000000100000001010101010101100;
		b = 32'b11010111010001110101100001100100;
		correct = 32'b01011000010010000110001000110001;
		#400 //-4.020834 * -219182450000000.0 = 881296200000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101101110110110101100100011100;
		b = 32'b00001111000011100101011000000101;
		correct = 32'b00111101011100111110101001000100;
		#400 //8.485618e+27 * 7.017707e-30 = 0.059549585
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011000100110101100010010110100;
		b = 32'b10101110000010001000011011001111;
		correct = 32'b01000111001001010001001111111111;
		#400 //-1361357000000000.0 * -3.1042554e-11 = 42259.996
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000110110001001101011010001110;
		b = 32'b01001000001101010101011101001001;
		correct = 32'b01001111100010110110111011001111;
		#400 //25195.277 * 185693.14 = 4678590000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010110000011001001100001001000;
		b = 32'b11011010010110111100010101011010;
		correct = 32'b10110000111100010110010101010000;
		#400 //1.1357161e-25 * -1.5465003e+16 = -1.7563853e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101100011000111000010000011001;
		b = 32'b00100101001001011111011111111010;
		correct = 32'b11010010000100111000000010000111;
		#400 //-1.1001999e+27 * 1.4395486e-16 = -158379130000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011010111101011011011000100010;
		b = 32'b10110001110110011011010111011011;
		correct = 32'b11001101010100001111010111101111;
		#400 //3.4580813e+16 * -6.336206e-09 = -219111150.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011111010010110111001011011011;
		b = 32'b01011111000111100001011101011011;
		correct = 32'b01111110111110110100011011100110;
		#400 //1.466002e+19 * 1.1391674e+19 = 1.6700218e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010100100100000010100011011111;
		b = 32'b11001000101011001101110010100100;
		correct = 32'b11011101110000101010111101101011;
		#400 //4953288000000.0 * -354021.12 = -1.7535686e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101100000100101010111100111010;
		b = 32'b00101011101110010000011011001111;
		correct = 32'b10011000010101000000100100001111;
		#400 //-2.0845118e-12 * 1.314693e-12 = -2.7404931e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010100010011000010001101001000;
		b = 32'b01000101001000000100111101010101;
		correct = 32'b10011001111111111010101010011111;
		#400 //-1.0306326e-26 * 2564.9583 = -2.6435295e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001111111101010110011101010101;
		b = 32'b00101100011100110001010111010111;
		correct = 32'b00111100111010010000011000000101;
		#400 //8234380000.0 * 3.45445e-12 = 0.028445253
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110101011111011011011011101100;
		b = 32'b10100011111110110100111010111011;
		correct = 32'b00011001111110010001000001100000;
		#400 //-9.451603e-07 * -2.7246818e-17 = 2.575261e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010111101100111110101011111000;
		b = 32'b01100011010001111011100101000011;
		correct = 32'b11111011100011000101110111011011;
		#400 //-395643530000000.0 * 3.6842516e+21 = -1.4576504e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111101000100000010011000111001;
		b = 32'b01000000010111001011010111001011;
		correct = 32'b00111101111110001000111001101101;
		#400 //0.035192702 * 3.4485958 = 0.121365406
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111111111110101000011000011011;
		b = 32'b10011011100111001111100010011101;
		correct = 32'b01111111111110101000011000011011;
		#400 //nan * -2.5968698e-22 = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111110011110011100110111110111;
		b = 32'b10010011100000101011000110110011;
		correct = 32'b01010010011111110000111111111011;
		#400 //-8.30118e+37 * -3.299184e-27 = 273871200000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010011000111111011001011100110;
		b = 32'b00110100110101001110011000010000;
		correct = 32'b10001000100001001100111110101011;
		#400 //-2.0156825e-27 * 3.965547e-07 = -7.9932835e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011101100010010011000100110111;
		b = 32'b11110110100011111011010100011010;
		correct = 32'b11010100100110100000011100010111;
		#400 //3.6314485e-21 * -1.4573665e+33 = -5292351300000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010100010010000011000110101101;
		b = 32'b11101000000001001111111010101001;
		correct = 32'b00111100110100000000000110000101;
		#400 //-1.01072164e-26 * -2.5122e+24 = 0.02539135
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100000010010001001101010001;
		b = 32'b00001011001110011010111110100110;
		correct = 32'b00001111110001101101101000000101;
		#400 //548.3018 * 3.5761847e-32 = 1.9608285e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101001111100010111110101100010;
		b = 32'b01011110000000111110101000000010;
		correct = 32'b01001000011110001101111111001111;
		#400 //1.07243004e-13 * 2.376353e+18 = 254847.23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010101011011100101011100000011;
		b = 32'b01111010101011001111110011010010;
		correct = 32'b11010000101000010000110111010111;
		#400 //-4.8132357e-26 * 4.4910143e+35 = -21616310000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000010100101110010101111101001;
		b = 32'b01011001111011110100110011000000;
		correct = 32'b00011101000011010100111101010001;
		#400 //2.221266e-37 * 8419613400000000.0 = 1.87022e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101101110000000000110001010010;
		b = 32'b01011100011011110101001100111011;
		correct = 32'b01001010101100111000100111110001;
		#400 //2.1833344e-11 * 2.6945613e+17 = 5883128.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111100100001001100100001011111;
		b = 32'b00001001111100100111010110000001;
		correct = 32'b11000110111110111000010010111001;
		#400 //-5.5155776e+36 * 5.836988e-33 = -32194.361
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101100101010011010101011100000;
		b = 32'b10100100111110110010100000111010;
		correct = 32'b11010010001001100111010100110011;
		#400 //1.6409232e+27 * -1.08922045e-16 = -178732710000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100101111000001110101110111001;
		b = 32'b11111001101010111011000000001011;
		correct = 32'b01100000000101101101100000100000;
		#400 //-3.9017538e-16 * -1.1143167e+35 = 4.347789e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011101100100111110010001011011;
		b = 32'b11000011101100101001110001001010;
		correct = 32'b00100001110011100101111000100010;
		#400 //-3.914669e-21 * -357.221 = 1.398402e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011000111010010111111101111000;
		b = 32'b00001000101010101111011110011001;
		correct = 32'b10100010000110111111000001111011;
		#400 //-2053869500000000.0 * 1.0289713e-33 = -2.1133726e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100110100010011111111100010000;
		b = 32'b10111101001010001100010110100111;
		correct = 32'b11100100001101011111001111011100;
		#400 //3.2583464e+23 * -0.04120412 = -1.342573e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101110111010000001011110010011;
		b = 32'b00010001011101000101110110010111;
		correct = 32'b11000000110111011000101101010010;
		#400 //-3.591451e+28 * 1.9277046e-28 = -6.923257
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111000011100101010011111100000;
		b = 32'b10100101010011110101111011010010;
		correct = 32'b11011110010001001000111110011111;
		#400 //1.9686574e+34 * -1.7986514e-16 = -3.5409285e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110010001111001110011111010;
		b = 32'b00100110010010001100111011101111;
		correct = 32'b10011101000111001001001111111110;
		#400 //-2.9744683e-06 * 6.9669386e-16 = -2.0722938e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011111001111100010001100011110;
		b = 32'b00101110001000000101110011101000;
		correct = 32'b00001101111011100011010111100111;
		#400 //4.0263113e-20 * 3.6462305e-11 = 1.4680859e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001010100101111000110010001100;
		b = 32'b01101110100001010110111001011011;
		correct = 32'b00111001100111011111101010110010;
		#400 //1.4593639e-32 * 2.064746e+28 = 0.00030132156
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110100001000100001001011000010;
		b = 32'b01100100010011101011010011001001;
		correct = 32'b11011001000000101101110110001101;
		#400 //-1.509425e-07 * 1.5252225e+22 = -2302209000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000000110111100100111000100100;
		b = 32'b10011101110010100001100111000100;
		correct = 32'b00011111001011111000000000001000;
		#400 //-6.9470387 * -5.3495596e-21 = 3.7163596e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101101101001100000101101010010;
		b = 32'b00101100010011011110111000110111;
		correct = 32'b11011010100001011001000110010011;
		#400 //-6.4235246e+27 * 2.9264488e-12 = -1.8798116e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010010000110001001000111001001;
		b = 32'b11000110011000110010110110101000;
		correct = 32'b00011001000001110110010001111011;
		#400 //-4.8142437e-28 * -14539.414 = 6.999628e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101100010100010110011101010010;
		b = 32'b11100110110001001001110111011001;
		correct = 32'b11010011101000001101010000111001;
		#400 //2.975804e-12 * -4.642478e+23 = -1381510500000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111100000010100010101100111001;
		b = 32'b10001101000001001111001100101100;
		correct = 32'b01001001100011111000001100010000;
		#400 //-2.8696545e+36 * -4.096835e-31 = 1175650.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010010011010011101100111110111;
		b = 32'b01111111110100111001100101111110;
		correct = 32'b01111111110100111001100101111110;
		#400 //-251096060000.0 * nan = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011000011110010111010111000;
		b = 32'b01010010101110000100011111101010;
		correct = 32'b11011110010011100010001110011010;
		#400 //-9383608.0 * 395740250000.0 = -3.7134713e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110101101011000110111110111100;
		b = 32'b11000001110111011110010011101101;
		correct = 32'b01111000000101010111011010101000;
		#400 //-4.3717837e+32 * -27.73678 = 1.212592e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111101001101100010100111101110;
		b = 32'b10011101001111010011101111101010;
		correct = 32'b11011011000001101010011110010111;
		#400 //1.5133575e+37 * -2.5044917e-21 = -3.7901914e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001110111110100100101110100100;
		b = 32'b01001011101101110000001010101101;
		correct = 32'b11011011001100101110111010110000;
		#400 //-2099630600.0 * 23987546.0 = -5.0364986e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010011101001001110011001001111;
		b = 32'b01111010010101101100010111010100;
		correct = 32'b11001110100010100101011111110100;
		#400 //-4.1626522e-27 * 2.7879099e+35 = -1160510000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000111100101100011111000011110;
		b = 32'b11101110110011111111100100101010;
		correct = 32'b10110110111101000001110011101011;
		#400 //2.2606e-34 * -3.218231e+28 = -7.275133e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000111010011010111010110101000;
		b = 32'b11000010110011011111010101101010;
		correct = 32'b10001010101001010100110000101110;
		#400 //1.5457062e-34 * -102.979324 = -1.5917578e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011011001111100010011101000001;
		b = 32'b11111010000111101000000010001001;
		correct = 32'b11010101111010110111011101100111;
		#400 //1.5729115e-22 * -2.0574748e+35 = -32362258000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010100101001101111111110110001;
		b = 32'b01001010001101010110010101111011;
		correct = 32'b00011111011011001010100111110111;
		#400 //1.6862569e-26 * 2971998.8 = 5.0115536e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100000010110000111101111101100;
		b = 32'b01000010001000000110001110100001;
		correct = 32'b10100011000001111010000110110100;
		#400 //-1.8336914e-19 * 40.097294 = -7.352607e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011101110011111110011000101000;
		b = 32'b01000100001101011011000110101010;
		correct = 32'b01100010100100111000111000000010;
		#400 //1.8725881e+18 * 726.776 = 1.360952e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111111111010111001110100000001;
		b = 32'b00111001101101010000000111101111;
		correct = 32'b10111010001001101001011111001001;
		#400 //-1.8407289 * 0.0003452445 = -0.0006355015
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011111011010000011000111111111;
		b = 32'b11111110011011100100100100111001;
		correct = 32'b01011110010110000010000011100101;
		#400 //-4.9169267e-20 * -7.9184114e+37 = 3.8934248e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010100101001011111100101010011;
		b = 32'b00110101000101100100011110001101;
		correct = 32'b01001010010000101101110011110100;
		#400 //5702820600000.0 * 5.5983475e-07 = 3192637.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101010011010110100111000101100;
		b = 32'b11001101101110010000111110010010;
		correct = 32'b01111000101010100001100111001110;
		#400 //-7.111668e+25 * -388100670.0 = 2.7600433e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010101011100000011101101111001;
		b = 32'b01101101011001101011010111011111;
		correct = 32'b01000011010110001000000000011010;
		#400 //4.851453e-26 * 4.4625888e+27 = 216.5004
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101101100010000010110011101010;
		b = 32'b01101101111000110010101101110001;
		correct = 32'b01011011111100011010110111011110;
		#400 //1.5481356e-11 * 8.788202e+27 = 1.3605328e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100101001100001111011000110111;
		b = 32'b01100100010000000011010001001010;
		correct = 32'b01001010000001001101110011001110;
		#400 //1.5348987e-16 * 1.4182171e+22 = 2176819.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000101011010001001010111010100;
		b = 32'b00111001000100101101010101010011;
		correct = 32'b00111111000001010110011101000011;
		#400 //3721.3643 * 0.00014003114 = 0.5211069
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110110000100101100000000101101;
		b = 32'b10111011101000010011010110110000;
		correct = 32'b11110010001110001101001101000110;
		#400 //7.441144e+32 * -0.00491973 = -3.660842e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000101110010010100011010000111;
		b = 32'b01000100011000111110001100000100;
		correct = 32'b01001010101100110010110000000110;
		#400 //6440.816 * 911.5471 = 5871107.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111001101001111101000000001110;
		b = 32'b10100101011011010011011000001111;
		correct = 32'b01011111100110110111111100001101;
		#400 //-1.0891668e+35 * -2.0574789e-16 = 2.2409377e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111111001000011011001011000100;
		b = 32'b00000001110011001010101101011010;
		correct = 32'b10000001100000010100011010101111;
		#400 //-0.631634 * 7.518364e-38 = -4.748854e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011111001000010110010101011101;
		b = 32'b01000011100000100000000100111100;
		correct = 32'b00100011001000111110110010000001;
		#400 //3.4176922e-20 * 260.00964 = 8.886329e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011111011011110010100110100011;
		b = 32'b10110110101001101010101111110000;
		correct = 32'b01010110100110111011010110100001;
		#400 //-1.7233485e+19 * -4.9672017e-06 = 85602200000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010100000000001101010011010011;
		b = 32'b11010110001101100001001001110100;
		correct = 32'b01101010101101110100000100101111;
		#400 //-2213305600000.0 * -50047593000000.0 = 1.1077062e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101000010111101111010010000010;
		b = 32'b01001110000101001001010101001000;
		correct = 32'b01110111000000010110011101011110;
		#400 //4.211503e+24 * 623202800.0 = 2.6246204e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101101001010011011001000000110;
		b = 32'b10100101001100011101000001111001;
		correct = 32'b01010010111010111011110010001110;
		#400 //-3.2823865e+27 * -1.5422936e-16 = 506240370000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000110011010110100100011110010;
		b = 32'b10101110011011101000010001100111;
		correct = 32'b00110101010110110011011110000001;
		#400 //-15058.236 * -5.423253e-11 = 8.1664626e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100011111100000011010011010111;
		b = 32'b10100100100100111110000110010011;
		correct = 32'b00001001000010101100001000000000;
		#400 //-2.604323e-17 * -6.4133225e-17 = 1.6702364e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111111000110110111010110001000;
		b = 32'b01110010101111000001010111000111;
		correct = 32'b11110010011001000110111100010011;
		#400 //-0.60726213 * 7.450817e+30 = -4.5245992e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111110100101000011111010010010;
		b = 32'b10000110001010001101101101100111;
		correct = 32'b01000101010000111001000000111010;
		#400 //-9.852531e+37 * -3.175848e-35 = 3129.0142
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101100111001100001101111111011;
		b = 32'b01010000101111000000110000111011;
		correct = 32'b01111110001010010000011110001011;
		#400 //2.2254806e+27 * 25239345000.0 = 5.6169674e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001110101000100011010010111100;
		b = 32'b00100010100110001010010010010111;
		correct = 32'b10110001110000010110111100110010;
		#400 //-1360682500.0 * 4.137395e-18 = -5.6296807e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111000000010001111000011110100;
		b = 32'b00010000010000111001101110010101;
		correct = 32'b01001000110100010100010110000111;
		#400 //1.1109992e+34 * 3.8576825e-29 = 428588.22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101011100100110011010100100001;
		b = 32'b11000001100100101111111011111001;
		correct = 32'b11101101101010010000110111010101;
		#400 //3.5592598e+26 * -18.374498 = -6.539961e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100111001010001011001111010000;
		b = 32'b01101011100111000111001100100110;
		correct = 32'b01010011010011100011001011101001;
		#400 //2.341216e-15 * 3.782724e+26 = 885617400000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111011110011111011100111111001;
		b = 32'b10110110010100000110111100000011;
		correct = 32'b01110010101010010010000100101110;
		#400 //-2.1571548e+36 * -3.1059033e-06 = 6.699914e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100101001110010100011110110100;
		b = 32'b10000011000000101101101000101010;
		correct = 32'b10101000101111010110100010011110;
		#400 //5.468503e+22 * -3.8454006e-37 = -2.1028586e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110001100110001110100010001010;
		b = 32'b01100110001110100100000100001000;
		correct = 32'b01011000010111100111111110011000;
		#400 //4.450219e-09 * 2.1988995e+23 = 978558400000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000001110110101110101001011000;
		b = 32'b01001010000010110010100100100100;
		correct = 32'b01001100011011100000000011011000;
		#400 //27.364426 * 2280009.0 = 62391136.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111101101011110101110010011101;
		b = 32'b00110011100110101111110101001101;
		correct = 32'b10110001110101000101011001110011;
		#400 //-0.085625865 * 7.217259e-08 = -6.17984e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001100101111010001110111111110;
		b = 32'b00111011001010000100100100001010;
		correct = 32'b01001000011110001010001101000111;
		#400 //99151860.0 * 0.00256783 = 254605.11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101101000110111100001101001011;
		b = 32'b01011101011010101000000011001110;
		correct = 32'b11001011000011101010111011100010;
		#400 //-8.854094e-12 * 1.0561083e+18 = -9350882.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111011100000100001000101001100;
		b = 32'b10110100010100110111111100100001;
		correct = 32'b00110000010101101110100110110010;
		#400 //-0.003969347 * -1.9697156e-07 = 7.818485e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010100110000101100111001111000;
		b = 32'b11000001110100110011111010000010;
		correct = 32'b11010111001000001011111110111110;
		#400 //6693501000000.0 * -26.405521 = -176745390000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101110101001110010000001111011;
		b = 32'b10011110111100111010000100101010;
		correct = 32'b01001110000111110000110100001100;
		#400 //-2.5861632e+28 * -2.5795282e-20 = 667108100.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100010001011101110110110000011;
		b = 32'b01001011011011011101110111011011;
		correct = 32'b00101110001000101000100101111011;
		#400 //2.3707135e-18 * 15588827.0 = 3.6956643e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101101110010011011000001001111;
		b = 32'b11101110111001010111110001000110;
		correct = 32'b11011101001101001100110010011111;
		#400 //2.2929351e-11 * -3.5511152e+28 = -8.1424767e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011100000011110101010001010001;
		b = 32'b00110111011111100011001001011111;
		correct = 32'b00010100000011100101000111011100;
		#400 //4.7423707e-22 * 1.5151308e-05 = 7.185312e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000010010100100000100111001011;
		b = 32'b10101001100000000000010011100100;
		correct = 32'b00101100010100100001000111010001;
		#400 //-52.509563 * -5.68519e-14 = 2.9852685e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000011101110000100010101101011;
		b = 32'b10011000100011100100101111110011;
		correct = 32'b00011100110011001101101001011001;
		#400 //-368.54233 * -3.678283e-24 = 1.3556029e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010111001100111000010011011001;
		b = 32'b00000011111101000101111000101000;
		correct = 32'b10011011101010110101110010100110;
		#400 //-197383160000000.0 * 1.4362648e-36 = -2.834945e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100001110001111011010100110100;
		b = 32'b10100011110101000000111001100011;
		correct = 32'b01000110001001010110110101001000;
		#400 //-4.604949e+20 * -2.2991179e-17 = 10587.32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000101111010011110101010110100;
		b = 32'b10101110100111110100111111101101;
		correct = 32'b00110101000100011001000111001110;
		#400 //-7485.338 * -7.2446805e-11 = 5.4228883e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010010010001011000000010001101;
		b = 32'b00000101001010110001010001000010;
		correct = 32'b00011000000000111111110001111111;
		#400 //212066320000.0 * 8.044102e-36 = 1.7058831e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111110001110100110101110010110;
		b = 32'b11100001000001011000111110010000;
		correct = 32'b01011111110000101000010011100000;
		#400 //-0.18205103 * -1.539851e+20 = 2.8033148e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011001100101010010111001000;
		b = 32'b10100010010111110111101101011000;
		correct = 32'b00101110000110111111010001111100;
		#400 //-11707848.0 * -3.0287433e-18 = 3.5460065e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000000100001011001111110100101;
		b = 32'b11011100110001101100111011010111;
		correct = 32'b00011101110011111000101011100001;
		#400 //-1.227139e-38 * -4.4767575e+17 = 5.493604e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101010100101001111011100011111;
		b = 32'b00000001101000101111111011001000;
		correct = 32'b00101100101111011011000101000110;
		#400 //9.004401e+25 * 5.9874995e-38 = 5.3913844e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100011001010011110111110011101;
		b = 32'b10001111111101110101011100000010;
		correct = 32'b00110011101001000010111111110010;
		#400 //-3.1347657e+21 * -2.4389595e-29 = 7.645566e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101100011111100100111101010101;
		b = 32'b00100011100000110000011000000000;
		correct = 32'b01010000100000100010100010001110;
		#400 //1.2297672e+27 * 1.420559e-17 = 17469567000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111000011010101111100100001110;
		b = 32'b00101111101010011111100001011001;
		correct = 32'b11101000100111000000001001011101;
		#400 //-1.9063264e+34 * 3.0917383e-10 = -5.893862e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000000010111101000111100101011;
		b = 32'b01110010110100010000111101010110;
		correct = 32'b11110011101101011100000000110111;
		#400 //-3.4774883 * 8.281716e+30 = -2.879957e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111100000110000101011111011111;
		b = 32'b10110011101100111100011011010111;
		correct = 32'b00110000010101011111011110001010;
		#400 //-0.009298294 * -8.371506e-08 = 7.784072e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110110000011011010001000111111;
		b = 32'b00100110110110001010100000111101;
		correct = 32'b11011101011011111011101111110011;
		#400 //-7.1816855e+32 * 1.5033612e-15 = -1.07966675e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111010101100100011100101000001;
		b = 32'b10111111011111000110100001110010;
		correct = 32'b11111010101011111011100100010011;
		#400 //4.6269504e+35 * -0.9859687 = -4.5620285e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111101000110011101111101000110;
		b = 32'b00111001000010011001010000100000;
		correct = 32'b10110110101001010110001100001010;
		#400 //-0.037566446 * 0.00013120519 = -4.928913e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100000010000001000110110101001;
		b = 32'b10001100010010110101111011100111;
		correct = 32'b10101101000110001111011110110111;
		#400 //5.5499727e+19 * -1.566711e-31 = -8.695203e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111111001010101001100111011111;
		b = 32'b00111111100100100011111000001100;
		correct = 32'b01111111010000101110101000110101;
		#400 //2.267677e+38 * 1.1425185 = 2.590863e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111010100010011111000011100001;
		b = 32'b11000001000011010001010100111011;
		correct = 32'b01111100000110000000101000111001;
		#400 //-3.5811514e+35 * -8.817683 = 3.157746e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000000101001100111011111101100;
		b = 32'b11111011101110110110101011000100;
		correct = 32'b01111100111100111011111000001101;
		#400 //-5.202139 * -1.94625e+36 = 1.01246626e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100101011000100111000000011010;
		b = 32'b11010100001001100110111110011001;
		correct = 32'b00111010000100110011011101100111;
		#400 //-1.9640357e-16 * -2859347500000.0 = 0.00056158606
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101001010011001110101101110001;
		b = 32'b10000011011110111110000010000011;
		correct = 32'b00101101010010011001111010001111;
		#400 //-1.5483294e+25 * -7.4019997e-37 = 1.1460734e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011010000010110110111011011010;
		b = 32'b01001110011011110110010011000011;
		correct = 32'b00101001000000100110001101011111;
		#400 //2.883407e-23 * 1004089540.0 = 2.895199e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011100001101101000000010101110;
		b = 32'b10010010010010001001010000110011;
		correct = 32'b10101111000011101111111000101111;
		#400 //2.0547972e+17 * -6.329154e-28 = -1.3005129e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100010110000001100010011000;
		b = 32'b11101110101110010100000110001100;
		correct = 32'b11110011100111000110000100011010;
		#400 //864.3843 * -2.8666984e+28 = -2.477929e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111111100001000010001111110101;
		b = 32'b11010001111000110100111101010001;
		correct = 32'b01010001111010101010100110100110;
		#400 //-1.0323473 * -122036036000.0 = 125983570000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010000001110001111000100001100;
		b = 32'b11100011100010011100101111000100;
		correct = 32'b00110100010001110001100001101000;
		#400 //-3.6473297e-29 * -5.0837736e+21 = 1.8542198e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110111010111000011111001100010;
		b = 32'b00001011100000110100101110010000;
		correct = 32'b11000011011000011110100111011101;
		#400 //-4.4670726e+33 * 5.057306e-32 = -225.91353
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011100110111111010000101101110;
		b = 32'b10110010001100010011100101110000;
		correct = 32'b01001111100110101101000011001010;
		#400 //-5.035713e+17 * -1.0315816e-08 = 5194749000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101111100010001101110110010001;
		b = 32'b11001110110010111110100000110001;
		correct = 32'b01111110110110100000011110101010;
		#400 //-8.471564e+28 * -1710495900.0 = 1.4490575e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101110110101111100000001110100;
		b = 32'b10010111111100001111110010001000;
		correct = 32'b00000111010010110001100101000001;
		#400 //-9.8112546e-11 * -1.5573384e-24 = 1.5279444e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101011010011111000111101111011;
		b = 32'b00100100110010001011010111000111;
		correct = 32'b10010000101000101011101101111010;
		#400 //-7.374029e-13 * 8.7044117e-17 = -6.4186587e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001110110111011000100100100001;
		b = 32'b01010011111111010101101011011010;
		correct = 32'b01100011010110110011111100100100;
		#400 //1858375800.0 * 2176301900000.0 = 4.0443867e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101111010101111011010010001111;
		b = 32'b10001001011001101011100111101101;
		correct = 32'b10111001010000100110100011100010;
		#400 //6.675756e+28 * -2.7772665e-33 = -0.00018540354
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101100111011100101110100110000;
		b = 32'b11110000110110000001011100011111;
		correct = 32'b11011110010010010011010000101000;
		#400 //6.7747127e-12 * -5.350137e+29 = -3.6245643e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100001111100101010010111010;
		b = 32'b01011011010100111001110011010000;
		correct = 32'b01100000000111010101010001101100;
		#400 //761.32385 * 5.9563637e+16 = 4.534722e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100000111000001011000110110010;
		b = 32'b00110011001110010001000011010111;
		correct = 32'b01010100101000100110111100110001;
		#400 //1.2952734e+20 * 4.3088985e-08 = 5581201500000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101010010110100100100100110100;
		b = 32'b01001010010010101011101011000010;
		correct = 32'b11110101001011001101110100000010;
		#400 //-6.597288e+25 * 3321520.5 = -2.1913028e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111100101000101100101111011101;
		b = 32'b11110010101011101000111110100001;
		correct = 32'b11101111110111100000001111001101;
		#400 //0.0198726 * -6.9150756e+30 = -1.3742053e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001100000000011000001001100011;
		b = 32'b00001101101110010101101000111111;
		correct = 32'b10011010001110111000100111000011;
		#400 //-33950092.0 * 1.1423231e-30 = -3.8781977e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001101011101101110010110101011;
		b = 32'b01010111001111000001100010111100;
		correct = 32'b00100101001101010110100010000100;
		#400 //7.6081055e-31 * 206814420000000.0 = 1.5734659e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100110000110110100010100110110;
		b = 32'b00011110100111111000110111110000;
		correct = 32'b10000101010000011000110000100110;
		#400 //-5.3870226e-16 * 1.6893484e-20 = -9.1005576e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111011001001110100111001000101;
		b = 32'b01001001000010111101000010010010;
		correct = 32'b11000100101101101011111110011101;
		#400 //-0.002552883 * 572681.1 = -1461.9879
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111011001100001100010000110100;
		b = 32'b10111011010101100011111111010101;
		correct = 32'b10110111000100111111000000010111;
		#400 //0.0026972415 * -0.0032691855 = -8.817783e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100100100100001001011000010010;
		b = 32'b10000110101101011001000010000110;
		correct = 32'b00101011110011010001011101110110;
		#400 //-2.1337159e+22 * -6.829699e-35 = 1.4572638e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100101110100111010010000100110;
		b = 32'b11001110101011100100110011011001;
		correct = 32'b00110101000100000001100100011010;
		#400 //-3.6713897e-16 * -1462135900.0 = 5.368071e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010111110111100110100001111100;
		b = 32'b10001110010011000000000111110100;
		correct = 32'b00100110101100010011110011110101;
		#400 //-489080680000000.0 * -2.5145882e-30 = 1.2298365e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111000100101101001010011001100;
		b = 32'b10110000111001010110100000011101;
		correct = 32'b11101010000001101111000001011000;
		#400 //2.4433203e+34 * -1.6691534e-09 = -4.0782763e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010101011000001101111101001111;
		b = 32'b01000110000100101001101101110000;
		correct = 32'b10011100000000001100011111100101;
		#400 //-4.54126e-26 * 9382.859 = -4.2610005e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001011101010101101101111110110;
		b = 32'b01011001110110100111110101011110;
		correct = 32'b10100110000100011101001011111100;
		#400 //-6.581258e-32 * 7687423500000000.0 = -5.059292e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100110111011010110000001000110;
		b = 32'b10110010100110001011001010111111;
		correct = 32'b11011010000011011001011011101000;
		#400 //5.604884e+23 * -1.7776413e-08 = -9963474000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101011110100100010000000111100;
		b = 32'b00111011010110001111010100010111;
		correct = 32'b00100111101100100001010001011110;
		#400 //1.4930344e-12 * 0.003310507 = 4.9427007e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110111111000111101100100110001;
		b = 32'b00001011011000001010000000101110;
		correct = 32'b11000011110001111110110010011100;
		#400 //-9.2426293e+33 * 4.3261337e-32 = -399.8485
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001110001001110011111010111101;
		b = 32'b01010000001100101101111000111111;
		correct = 32'b10011110111010011011010110100010;
		#400 //-2.0614547e-30 * 12003638000.0 = -2.4744956e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101011010000100000011001111100;
		b = 32'b00111001001100110001010111001100;
		correct = 32'b01100101000001111011101100001110;
		#400 //2.3456223e+26 * 0.0001707889 = 4.0060627e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111011110010100111101011111000;
		b = 32'b00110001110111100011011010110110;
		correct = 32'b01101110001011111100000111101001;
		#400 //2.1026761e+36 * 6.4672703e-09 = 1.3598575e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111101001011111101000101011;
		b = 32'b00111011101101001001101111001101;
		correct = 32'b10110011111010100011000111010011;
		#400 //-1.9786026e-05 * 0.005511737 = -1.0905537e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110110101110001010110111010111;
		b = 32'b10100101001111001011010100111010;
		correct = 32'b10011100100010000010001001100111;
		#400 //5.503865e-06 * -1.6367803e-16 = -9.008618e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001111100000100011101000011010;
		b = 32'b11100001000001110101101111101101;
		correct = 32'b10110001000010011011011011001110;
		#400 //1.284137e-29 * -1.560584e+20 = -2.0040036e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010100111001111001101010000010;
		b = 32'b10110000011001111100000101010110;
		correct = 32'b00000101110100011010101101010101;
		#400 //-2.3385982e-26 * -8.431206e-10 = 1.9717203e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100111101000000000011111011010;
		b = 32'b00011101000011110100111010001001;
		correct = 32'b00000101001100110010101011110110;
		#400 //4.4417434e-15 * 1.8966494e-21 = 8.42443e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110110100001110010100011011010;
		b = 32'b00000100011011100010000100010100;
		correct = 32'b00111011011110110111001011100011;
		#400 //1.370681e+33 * 2.7991954e-36 = 0.0038368038
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110100111100101000011101110;
		b = 32'b01100101000110011000010011101110;
		correct = 32'b11011100001111011110000100100110;
		#400 //-4.7181884e-06 * 4.5310887e+22 = -2.137853e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010011110101000101110101011101;
		b = 32'b01010000111010110111010100110001;
		correct = 32'b10100101010000110101001011101100;
		#400 //-5.3608387e-27 * 31602608000.0 = -1.6941649e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111001001110101011010110110101;
		b = 32'b00100010110110100001000010011100;
		correct = 32'b11011100100111110000101011011001;
		#400 //-6.059079e+34 * 5.9106604e-18 = -3.581316e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110001001001100111001000100111;
		b = 32'b00011010000111001001000011101001;
		correct = 32'b10001011110010111001011110001111;
		#400 //-2.4221067e-09 * 3.23771e-23 = -7.8420796e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001111111110110111100110110101;
		b = 32'b11011110001010000110101101011111;
		correct = 32'b01101110101001010111000101011000;
		#400 //-8438115000.0 * -3.0339745e+18 = 2.5601025e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001110100010000000001110001001;
		b = 32'b10100001101010001100001101101101;
		correct = 32'b10110000101100110101010001001101;
		#400 //1140966500.0 * -1.1435852e-18 = -1.3047924e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110010001001011110101000011100;
		b = 32'b11000111001011011000001000110001;
		correct = 32'b11111001111000001110011100101011;
		#400 //3.286275e+30 * -44418.19 = -1.4597039e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011001001110110000000110000110;
		b = 32'b00110001100001010111000010001001;
		correct = 32'b11001011010000101111001111111111;
		#400 //-3289843500000000.0 * 3.883603e-09 = -12776447.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111010100001011001111111100101;
		b = 32'b10100101011100100011010011000111;
		correct = 32'b11100000011111001101100101100110;
		#400 //3.4690926e+35 * -2.1008036e-16 = -7.2878824e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011101100110010111001000111110;
		b = 32'b01110011000011111011010111000111;
		correct = 32'b01010001001011000100011110001011;
		#400 //4.0616886e-21 * 1.1385885e+31 = 46245917000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110100001010111001001101100;
		b = 32'b00010010010110101000101100110000;
		correct = 32'b10001001011000111101011111111100;
		#400 //-3.9770293e-06 * 6.8960233e-28 = -2.7425686e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111010101111100100010101111011;
		b = 32'b10011010110101100111011110100001;
		correct = 32'b11010110000111110110011011111111;
		#400 //4.939728e+35 * -8.8701596e-23 = -43816180000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001101011010101110111111111010;
		b = 32'b11011101110100010110111100100010;
		correct = 32'b01101011110000000011001111101000;
		#400 //-246349730.0 * -1.8864148e+18 = 4.6471776e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010110110111101001100001100000;
		b = 32'b11101111110000110011101100111111;
		correct = 32'b11000111001010011100000110010101;
		#400 //3.5962197e-25 * -1.208424e+29 = -43457.582
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101011100100000001110100101100;
		b = 32'b01101100100111100001101111110110;
		correct = 32'b01011000101100100000001101111101;
		#400 //1.0239912e-12 * 1.5291386e+27 = 1565824400000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110101000010101011011000000000;
		b = 32'b10001100000110111110000101001101;
		correct = 32'b10000001101010001110110010001011;
		#400 //5.167385e-07 * -1.2008565e-31 = -6.2052876e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000011011110111001001111000001;
		b = 32'b01011111100110111011000111111011;
		correct = 32'b10100011100110010000000101011110;
		#400 //-7.3931884e-37 * 2.2438048e+19 = -1.6588872e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011011110110110000010010100001;
		b = 32'b10101000101000110010011001001111;
		correct = 32'b10000101000010111001010010111001;
		#400 //3.6233502e-22 * -1.8113249e-14 = -6.5630646e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001111111011101110110000000010;
		b = 32'b01010001110001010001110111100111;
		correct = 32'b01100010001101111111011110000110;
		#400 //8016889000.0 * 105826280000.0 = 8.483975e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000000101001011001111101101110;
		b = 32'b01111100000101111011010001111001;
		correct = 32'b01111101010001000100101110011001;
		#400 //5.1757116 * 3.150789e+36 = 1.6307576e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010111101100011000110101100001;
		b = 32'b00011111000001000100011110110011;
		correct = 32'b10110111001101110111110101000001;
		#400 //-390441550000000.0 * 2.8011395e-20 = -1.0936813e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010001100010010110001010001101;
		b = 32'b10111001111001010011100010000111;
		correct = 32'b01001011111101100000011011111100;
		#400 //-73757990000.0 * -0.000437204 = 32247288.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111010100110010010111011111;
		b = 32'b10011000100110110111011110101010;
		correct = 32'b10100000100000000011101010100001;
		#400 //54053.87 * -4.018739e-24 = -2.172284e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100111110111010011000000000110;
		b = 32'b11000101000101100000110111001001;
		correct = 32'b01101101100000011010011000001101;
		#400 //-2.0890577e+24 * -2400.8616 = 5.0155387e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101101110001000101001100100011;
		b = 32'b11011010010000010111110011001101;
		correct = 32'b11001000100101000110001001100011;
		#400 //2.231954e-11 * -1.3615473e+16 = -303891.1
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010100010011101000001100011001;
		b = 32'b00111010011001111010010000111000;
		correct = 32'b01001111001110101101110011000101;
		#400 //3547850900000.0 * 0.0008836421 = 3135030500.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111101111001110101110001101100;
		b = 32'b10111010010100001010011111101110;
		correct = 32'b11111000101111001001001011011100;
		#400 //3.8441444e+37 * -0.0007959594 = -3.0597827e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010100111101100111010001011101;
		b = 32'b00010101111000011001010110001010;
		correct = 32'b00101011010110010010110000111100;
		#400 //8468113700000.0 * 9.111271e-26 = 7.7155274e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000111001101111010011100010111;
		b = 32'b01111101110110110111111111001110;
		correct = 32'b01000101100111010111011110100000;
		#400 //1.3816493e-34 * 3.6470566e+37 = 5038.953
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101110001001000010010100100010;
		b = 32'b00100000010000001101101100010100;
		correct = 32'b01001110111101110101000010100100;
		#400 //1.2700108e+28 * 1.633552e-19 = 2074628600.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101011101111011011110111011100;
		b = 32'b11111110110011001101101101010011;
		correct = 32'b01101011000101111101010111011010;
		#400 //-1.3481954e-12 * -1.3615065e+38 = 1.8355768e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001001110100011110010001101111;
		b = 32'b10111101110101001000001101011110;
		correct = 32'b11001000001011100011110011100001;
		#400 //1719437.9 * -0.10376619 = -178419.52
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011110101010110111000111111011;
		b = 32'b10110001111010000111010000011101;
		correct = 32'b11010001000110111010110100001111;
		#400 //6.1769656e+18 * -6.765289e-09 = -41788960000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000000011001111001110011100101;
		b = 32'b01100011010110001011100010110110;
		correct = 32'b01100100010001000001001101111111;
		#400 //3.618951 * 3.9978065e+21 = 1.4467867e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110000100010111010010100011110;
		b = 32'b11101100100010110100001010111101;
		correct = 32'b11011101100101111110111000011110;
		#400 //1.016051e-09 * -1.3468468e+27 = -1.3684651e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111100100011001101001110001;
		b = 32'b10100011101110100010011000110111;
		correct = 32'b00011011110100111011111111100101;
		#400 //-1.7357264e-05 * -2.0182345e-17 = 3.503103e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000011010001100110011111101001;
		b = 32'b01000001111110111011010111100101;
		correct = 32'b00000101110000110001010011011010;
		#400 //5.8306253e-37 * 31.463816 = 1.8345372e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101010000101001011100011110000;
		b = 32'b10101010000100111100110100011101;
		correct = 32'b10010100101010111011101010110110;
		#400 //1.3209204e-13 * -1.3127386e-13 = -1.7340232e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010110111100100000111110001;
		b = 32'b10101010001100101110011001101000;
		correct = 32'b00100101100110110101000111100011;
		#400 //-0.0016956908 * -1.5889514e-13 = 2.6943702e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111011111010010110101100111010;
		b = 32'b00101100011101011010101001001000;
		correct = 32'b01101000110111111111111011100001;
		#400 //2.42396e+36 * 3.491112e-12 = 8.4623153e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010100110100100010110110101111;
		b = 32'b00111110101010100101100001001011;
		correct = 32'b00010100000010111101101011010011;
		#400 //2.12226e-26 * 0.33270487 = 7.060862e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111001011001010011000001000101;
		b = 32'b10010100111110110111111010110000;
		correct = 32'b10001110111000010010011110111111;
		#400 //0.00021857124 * -2.5394493e-26 = -5.5505056e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111100001100010000111110110001;
		b = 32'b01101001111101110011100010001001;
		correct = 32'b11100110101010101111110100111110;
		#400 //-0.010806964 * 3.7358957e+25 = -4.037369e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011010010000100010100101100110;
		b = 32'b11000110101011111111100110110011;
		correct = 32'b00100001100001010111011110101111;
		#400 //-4.01517e-23 * -22524.85 = 9.044111e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110111010011100100001101101111;
		b = 32'b00101110000110111101001111100110;
		correct = 32'b00100101111110110001101100011110;
		#400 //1.2294257e-05 * 3.5431123e-11 = 4.3559935e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111111001010000110110000100100;
		b = 32'b10010010111001010010001001101111;
		correct = 32'b00010010100101101011111101100100;
		#400 //-0.6579001 * -1.446042e-27 = 9.513512e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010100001100001110110010110010;
		b = 32'b10001101100011101000101110001010;
		correct = 32'b10100010010001010000011101110101;
		#400 //3039541300000.0 * -8.7850185e-31 = -2.6702426e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011110010100100010101111100100;
		b = 32'b00110010010111101100100011101000;
		correct = 32'b01010001001101101110011100000000;
		#400 //3.7861122e+18 * 1.29677815e-08 = 49097474000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110000100100101011000011101100;
		b = 32'b00110100000101111001100101111011;
		correct = 32'b00100101001011011011110010011011;
		#400 //1.0673182e-09 * 1.4118807e-07 = 1.506926e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010111000001100101001011010110;
		b = 32'b11100110010010000000111110001101;
		correct = 32'b10111101110100011111000111000000;
		#400 //4.340229e-25 * -2.3619004e+23 = -0.10251188
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111010000000001001101111000001;
		b = 32'b00001110000000010011110111010011;
		correct = 32'b00001000100000011101101100010111;
		#400 //0.00049060216 * 1.5930245e-30 = 7.815413e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001010001110011111011010110000;
		b = 32'b11000110001100001011110110101001;
		correct = 32'b10010001000000000110001101011111;
		#400 //8.953823e-33 * -11311.415 = -1.0128041e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011100011110000101111100101011;
		b = 32'b10010010111100110000110011110111;
		correct = 32'b10101111111010111100111011101010;
		#400 //2.7964173e+17 * -1.5338652e-27 = -4.2893272e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011111110100100110111001110001;
		b = 32'b01011011000011000011101110011000;
		correct = 32'b00111011011001101000101011000100;
		#400 //8.912117e-20 * 3.947202e+16 = 0.0035177926
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101000011011011011111110011110;
		b = 32'b01000001010000101110000101000000;
		correct = 32'b01101010001101001111110001100111;
		#400 //4.4909423e+24 * 12.179993 = 5.4699646e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010001111010010100100011100001;
		b = 32'b01010110111000001111011010100011;
		correct = 32'b01101001010011010000000010000101;
		#400 //125243760000.0 * 123674950000000.0 = 1.5489515e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110011001100111100100010011011;
		b = 32'b01010000100000100000010111001110;
		correct = 32'b01000100001101101001111111100101;
		#400 //4.1859135e-08 * 17451348000.0 = 730.49835
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110100100011010001110111110010;
		b = 32'b00111111100011010110111010011110;
		correct = 32'b11110100100110111110110011110001;
		#400 //-8.944351e+31 * 1.1049383 = -9.882956e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110100010000000000100011101100;
		b = 32'b00111000100111000011010000010101;
		correct = 32'b01101101011010100101100100000011;
		#400 //6.0858274e+31 * 7.448361e-05 = 4.5329438e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000000111001111110001001010100;
		b = 32'b11011000010000110101110011111101;
		correct = 32'b10011001101100001111010110100000;
		#400 //2.1295191e-38 * -859216600000000.0 = -1.829718e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111101111111001000010010010000;
		b = 32'b00111111010101011100111010100110;
		correct = 32'b10111101110100101110011000100010;
		#400 //-0.12329972 * 0.83518445 = -0.102978006
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010001010011110100001010111011;
		b = 32'b01000110001101001101100010010101;
		correct = 32'b01011000000100100110101001000100;
		#400 //55636110000.0 * 11574.1455 = 643940400000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000010001110010100010010111110;
		b = 32'b10011101101101110000011000011001;
		correct = 32'b10100000100001000111010010001110;
		#400 //46.31713 * -4.8446e-21 = -2.24388e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011110100110001100110101010101;
		b = 32'b01010110101101101110000110011001;
		correct = 32'b01110101110110100101000101000100;
		#400 //5.505275e+18 * 100540025000000.0 = 5.5350048e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010100010001111101000010000010;
		b = 32'b11000001101110000010111011110010;
		correct = 32'b10010110100011111100001010000010;
		#400 //1.00880534e-26 * -23.022923 = -2.3225648e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000110110111011111101100101110;
		b = 32'b00001110111001001110110110111101;
		correct = 32'b00010110010001101000000111011010;
		#400 //28413.59 * 5.6435273e-30 = 1.6035287e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110000010000101001001011101001;
		b = 32'b10100001110001100111100010110100;
		correct = 32'b10010010100101101101100101011110;
		#400 //7.078556e-10 * -1.3448952e-18 = -9.519916e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100110100000111010001101011101;
		b = 32'b11101101001001111011000111000101;
		correct = 32'b11010100001011000111010111110110;
		#400 //9.134231e-16 * -3.2436817e+27 = -2962853700000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110100100111001110011110111111;
		b = 32'b01011011010001010110010111000011;
		correct = 32'b01010000011100011111100101101010;
		#400 //2.9225882e-07 * 5.556246e+16 = 16238619000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100111010110001001101000000010;
		b = 32'b10100011110111011110110110111000;
		correct = 32'b00001011101110111100011000010110;
		#400 //-3.005951e-15 * -2.4061546e-17 = 7.2327827e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001101000110010001111100101010;
		b = 32'b11100011011001100100111011000000;
		correct = 32'b00110001000010011100000100011010;
		#400 //-4.7184277e-31 * -4.2484257e+21 = 2.004589e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001001010100010111101111001011;
		b = 32'b00111101111100011001101000100110;
		correct = 32'b11000111110001011011001110101110;
		#400 //-858044.7 * 0.117969796 = -101223.36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001110110001101000001100000011;
		b = 32'b00100111010011110001110011010010;
		correct = 32'b00110110101000001001101001001001;
		#400 //1665237400.0 * 2.8742644e-15 = 4.7863327e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100011111101000100101111011010;
		b = 32'b00100010001010111010101001011111;
		correct = 32'b11000110101000111101000101000000;
		#400 //-9.0129425e+21 * 2.3265015e-18 = -20968.625
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100000111100010111001110011001;
		b = 32'b00111101001110110111100011110011;
		correct = 32'b00011110101100001101000110000100;
		#400 //4.0903484e-19 * 0.045769643 = 1.8721378e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110110011000011111000101111011;
		b = 32'b10110110111010100011000111010000;
		correct = 32'b11101101110011101011001010110001;
		#400 //1.14566855e+33 * -6.9795424e-06 = -7.996242e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000111110111001010111111100001;
		b = 32'b10000101110000111011001101000100;
		correct = 32'b00001110001010001011010010000010;
		#400 //-112991.76 * -1.8403564e-35 = 2.079451e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100111000010000100000011000101;
		b = 32'b00110011100010000000100111100100;
		correct = 32'b00011011000100001100111101011001;
		#400 //1.8908903e-15 * 6.3347926e-08 = 1.1978398e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111010000110010110101110100001;
		b = 32'b01000100000000001010001101110010;
		correct = 32'b00111110100110100010111110001001;
		#400 //0.0005852525 * 514.55383 = 0.3011439
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111001100010011011000101010110;
		b = 32'b10111011100100001000000100101011;
		correct = 32'b11110101100110110111001001110100;
		#400 //8.936768e+34 * -0.0044099293 = -3.9410517e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010110101001100010111110100001;
		b = 32'b11011001001110111010101010011111;
		correct = 32'b01110000011100111010011100011011;
		#400 //-91361750000000.0 * -3301463800000000.0 = 3.016275e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010000101011111011000000110101;
		b = 32'b01010101111110101111010010101100;
		correct = 32'b00100111001011000011100111111110;
		#400 //6.929682e-29 * 34491096000000.0 = 2.3901233e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010011111011100000100111100110;
		b = 32'b01100001110000000000101101011000;
		correct = 32'b10110110001100101001000111111001;
		#400 //-6.0089407e-27 * 4.4282403e+20 = -2.6609034e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010100011100001101001000011000;
		b = 32'b11010011111011011001111010001000;
		correct = 32'b10101000110111111000011110100010;
		#400 //1.2158337e-26 * -2041133900000.0 = -2.4816795e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011011100100100010001001101011;
		b = 32'b00000110100101011000100111110011;
		correct = 32'b00100010101010101011100110001111;
		#400 //8.226638e+16 * 5.625027e-35 = 4.627506e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000101110111001100011100011000;
		b = 32'b01001100011101111010011101111111;
		correct = 32'b01010010110101011001010010001100;
		#400 //7064.8867 * 64921084.0 = 458660120000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010111000110101011011110101011;
		b = 32'b11011010010110111101010010110010;
		correct = 32'b11110010000001001101101110101011;
		#400 //170113640000000.0 * -1.546922e+16 = -2.6315253e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111100001110101111001000100000;
		b = 32'b01001000000000010000011010110111;
		correct = 32'b01000100101111000111000111010011;
		#400 //0.011410266 * 132122.86 = 1507.557
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100001001000101010001000001110;
		b = 32'b01000011101010100111110011110000;
		correct = 32'b01100101010110001001110111111001;
		#400 //1.8750311e+20 * 340.97607 = 6.3934078e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111101011110001111110001010100;
		b = 32'b01100111001011011000110010100001;
		correct = 32'b01100101001010001100101101001011;
		#400 //0.060787514 * 8.1956355e+23 = 4.981923e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010011111010010101000001010101;
		b = 32'b10111111010111101110110100101010;
		correct = 32'b10010011110010110010101111001111;
		#400 //5.8896683e-27 * -0.87080634 = -5.1287603e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101001001101010100111001010111;
		b = 32'b01001100000111111110100111001100;
		correct = 32'b11110101111000101000001001111010;
		#400 //-1.3699095e+25 * 41920304.0 = -5.7427025e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001011010101011111101111110111;
		b = 32'b11100110111000101010111110001101;
		correct = 32'b10110010101111010111101100101101;
		#400 //4.1211865e-32 * -5.352466e+23 = -2.205851e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011000000011001111111000000100;
		b = 32'b01011010000010010000101000001100;
		correct = 32'b01110010100101101111001011110001;
		#400 //620090500000000.0 * 9643280000000000.0 = 5.9797056e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110101010011101101111111111010;
		b = 32'b00001100001110010111101000101111;
		correct = 32'b11000010000101011110001010011000;
		#400 //-2.622451e+32 * 1.428865e-31 = -37.471283
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110100100101111011100010001011;
		b = 32'b01000111110001100111010101000110;
		correct = 32'b11111100111010110011110001111001;
		#400 //-9.616453e+31 * 101610.55 = -9.7713303e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001010000011100010101000011010;
		b = 32'b11001101110010011110101011111111;
		correct = 32'b00011000011000000100001100011101;
		#400 //-6.84497e-33 * -423452640.0 = 2.8985205e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110110110000011111100011000100;
		b = 32'b11110111101000111000010111001110;
		correct = 32'b11101110111101111100110110001110;
		#400 //5.7808084e-06 * -6.633268e+33 = -3.834565e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000011001010110011110001000100;
		b = 32'b01100001100011001101011000110111;
		correct = 32'b11100101001111000110100001111101;
		#400 //-171.23541 * 3.247475e+20 = -5.5608273e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011111110100000011010110011101;
		b = 32'b11111000001111101000110101101110;
		correct = 32'b11011000100110101111101011010010;
		#400 //8.818012e-20 * -1.5459452e+34 = -1363216400000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011011010010001101010001000001;
		b = 32'b01001001111011111000011111101100;
		correct = 32'b00100101101110111110100011001010;
		#400 //1.6612195e-22 * 1962237.5 = 3.2597073e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010100011101000011111101111110;
		b = 32'b01100010101110100101000110000001;
		correct = 32'b11110111101100011100001111100101;
		#400 //-4196149000000.0 * 1.7184837e+21 = -7.211014e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100110100111101001101001110101;
		b = 32'b10011111111001111001010001011000;
		correct = 32'b11000111000011110111100101000111;
		#400 //3.7449157e+23 * -9.807772e-20 = -36729.277
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011101111110011110100011011111;
		b = 32'b00111111001010000111010111001101;
		correct = 32'b01011101101001000111001111010010;
		#400 //2.250986e+18 * 0.6580475 = 1.4812557e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001111000101001001001110101011;
		b = 32'b11110011111001101100110011010011;
		correct = 32'b01000011100001011111001110001100;
		#400 //-7.325403e-30 * -3.6571735e+31 = 267.9027
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011000001101011001010100000111;
		b = 32'b11000100010111010111011000101001;
		correct = 32'b01011101000111010001010101110111;
		#400 //-798606700000000.0 * -885.84625 = 7.0744276e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001100101110111000011000110110;
		b = 32'b10111110111111100010110101101101;
		correct = 32'b01001100001110100011000001110000;
		#400 //-98316720.0 * -0.49644032 = 48808384.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011101001111001010010001011010;
		b = 32'b10010001010101000100000000001111;
		correct = 32'b10101111000111000110011101001111;
		#400 //8.49568e+17 * -1.6743591e-28 = -1.422482e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110001010110000001111000000110;
		b = 32'b10000001000110001100010100010111;
		correct = 32'b00110011000000001111100000110110;
		#400 //-1.0701609e+30 * -2.8059396e-38 = 3.002807e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101000011001010011001000101110;
		b = 32'b01101000100010001000111001011100;
		correct = 32'b01010001011101001000010000111001;
		#400 //1.2722935e-14 * 5.158943e+24 = 65636897000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100000100100100101011101010110;
		b = 32'b00001100111001011111110101100110;
		correct = 32'b00101110000000110111100011111011;
		#400 //8.435993e+19 * 3.5435545e-31 = 2.9893404e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001001010011101010100100110000;
		b = 32'b00111100101001011111011001000110;
		correct = 32'b00000110100001011111100111011011;
		#400 //2.48759e-33 * 0.020259034 = 5.039617e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010111000010010111100001000111;
		b = 32'b11101001110100011011011111100001;
		correct = 32'b01000001011000010011101111100000;
		#400 //-4.44189e-25 * -3.169173e+25 = 14.077118
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000111110111010100111100011111;
		b = 32'b11111110100110001101010101011010;
		correct = 32'b01000111000001000001111101101011;
		#400 //-3.3298887e-34 * -1.0157522e+38 = 33823.418
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111110110111000001111010101001;
		b = 32'b00100100001110010110111100100101;
		correct = 32'b01100011100111110111000110111001;
		#400 //1.4629468e+38 * 4.0209623e-17 = 5.882454e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100001100010100101100111010;
		b = 32'b00000001101011110100011100100101;
		correct = 32'b00000110011100101100011101100100;
		#400 //709.1754 * 6.4386935e-38 = 4.566163e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111100010110110010000101110101;
		b = 32'b11111100101001010000100011110001;
		correct = 32'b01111001100011010100010000111000;
		#400 //-0.013374676 * -6.8552827e+36 = 9.168719e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001100111100011101111011001011;
		b = 32'b01111101110011110110001110001010;
		correct = 32'b11001011010000111111000100110010;
		#400 //-3.7266018e-31 * 3.445838e+37 = -12841266.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011110111100000100011101100011;
		b = 32'b01010111000101010011000000110011;
		correct = 32'b10110110100011000000011011001010;
		#400 //-2.5440513e-20 * 164034250000000.0 = -4.1731155e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010101001111101010010100100000;
		b = 32'b01111110010100011011001100110000;
		correct = 32'b11010100000111000010101001000000;
		#400 //-3.8500455e-26 * 6.968476e+37 = -2682895000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001100111101110110000111111010;
		b = 32'b00100111110101101111111011110000;
		correct = 32'b10110101010011111100001001000010;
		#400 //-129699790.0 * 5.9673336e-15 = -7.739619e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010101111110100100101111010011;
		b = 32'b01010011111110001010111001010011;
		correct = 32'b10101010011100110010001111100101;
		#400 //-1.01093825e-25 * 2136153100000.0 = -2.1595189e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001001111010011010010010000011;
		b = 32'b10110111010010101101011101110000;
		correct = 32'b01000001101110010010000001101111;
		#400 //-1914000.4 * -1.2090299e-05 = 23.140837
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101000111001010100011100001011;
		b = 32'b01100100101011100011110100101010;
		correct = 32'b11001110000111000000110100010001;
		#400 //-2.5454917e-14 * 2.5713126e+22 = -654525500.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110111011111111100101000000011;
		b = 32'b00101100110100110011011011010110;
		correct = 32'b01100100110100110000101001001011;
		#400 //5.1880195e+33 * 6.0030687e-12 = 3.1144037e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000101000011101111000000001010;
		b = 32'b00111100000000111111110000111101;
		correct = 32'b00000001100100110110001101010111;
		#400 //6.720896e-36 * 0.008055744 = 5.414182e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001011100100001110000001010100;
		b = 32'b11010001100110110111100111010100;
		correct = 32'b00011101101011111111100110001010;
		#400 //-5.5804314e-32 * -83470480000.0 = 4.658013e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000110100011111000000011011;
		b = 32'b10011111101111110000111101111001;
		correct = 32'b00010001000111001010111011010100;
		#400 //-1.5274993e-09 * -8.0917244e-20 = 1.2360103e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110011100110011101110001000101;
		b = 32'b01010000001001010111111101101000;
		correct = 32'b11000100010001101110111100010111;
		#400 //-7.1646845e-08 * 11106361000.0 = -795.7358
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110010011111001110001110001100;
		b = 32'b00110000001110101010000011011110;
		correct = 32'b11100011001110000101110000111101;
		#400 //-5.0089798e+30 * 6.789501e-10 = -3.4008474e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010000101011001100111101001100;
		b = 32'b00111010111001000001000110111011;
		correct = 32'b11001100000110011111010010011000;
		#400 //-23194132000.0 * 0.0017400304 = -40358496.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001010110011001110100100000010;
		b = 32'b11111110100100110100001110111110;
		correct = 32'b01001001111010111100000000001010;
		#400 //-1.9732133e-32 * -9.787413e+37 = 1931265.2
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000001110011000000001111000001;
		b = 32'b01111001111000000111000000011101;
		correct = 32'b01111100001100101101110010100010;
		#400 //25.501833 * 1.4566855e+35 = 3.7148152e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111111011011010011010001001100;
		b = 32'b10101110000101001101000010100000;
		correct = 32'b01101110000010011110001110001011;
		#400 //-3.1529858e+38 * -3.38366e-11 = 1.0668632e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011101010111000010111110000110;
		b = 32'b11011101101011100110100010111000;
		correct = 32'b11111011100101100000001001011111;
		#400 //9.9162796e+17 * -1.5709371e+18 = -1.5577852e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110000111000000011101111001100;
		b = 32'b01000100011011011110000010000001;
		correct = 32'b00110101110100000101110000000001;
		#400 //1.631514e-09 * 951.5079 = 1.5523984e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011100001011011001110111010000;
		b = 32'b11101010110001111100110111110010;
		correct = 32'b01000111100001111000000101011000;
		#400 //-5.7444866e-22 * -1.2077439e+26 = 69378.69
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111111100111010000111111100111;
		b = 32'b10000011101000100111110100010110;
		correct = 32'b00000011110001110110000110011101;
		#400 //-1.2270478 * -9.550223e-37 = 1.171858e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010000111100001011100011101001;
		b = 32'b00111110110111101001010111101111;
		correct = 32'b01010000010100010100110101010110;
		#400 //32309200000.0 * 0.43473765 = 14046026000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101101111110110010000011000100;
		b = 32'b00101011101101010010100001000011;
		correct = 32'b00011010001100011011010110101001;
		#400 //2.8549947e-11 * 1.2871998e-12 = 3.6749486e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100101101100010000100000010100;
		b = 32'b00110000000101111001001010011101;
		correct = 32'b10010110010100011010001001001110;
		#400 //-3.071008e-16 * 5.514183e-10 = -1.69341e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010011110010011101110110000001;
		b = 32'b10110001001000001011100010010011;
		correct = 32'b00000101011111010111011111110111;
		#400 //-5.0957953e-27 * -2.3387983e-09 = 1.1918037e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011101011001101101111010000011;
		b = 32'b01000010001111001001000101101111;
		correct = 32'b01100000001010100000111010010000;
		#400 //1.0397424e+18 * 47.142025 = 4.901556e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001000111111010011000100010110;
		b = 32'b00111100000111000011111011010010;
		correct = 32'b01000101100110101000100000001011;
		#400 //518536.7 * 0.009536462 = 4945.0054
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100011010000000011000000011011;
		b = 32'b10011111110111001100110011110111;
		correct = 32'b10000011101001011100001100110111;
		#400 //1.04185276e-17 * -9.351271e-20 = -9.7426475e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010010111000100110010000010001;
		b = 32'b11000000101001100101011011011100;
		correct = 32'b01010100000100110001100110110011;
		#400 //-486170720000.0 * -5.198103 = 2527165400000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100010000110110111111000100101;
		b = 32'b11101110011110101001111011101010;
		correct = 32'b01010001000110000011100110110110;
		#400 //-2.1073197e-18 * -1.9390842e+28 = 40862704000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110111011111001001010101010110;
		b = 32'b10111010000100000100110001100101;
		correct = 32'b01110010000011100101111101100000;
		#400 //-5.1229988e+33 * -0.0005504548 = 2.819979e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101001001001100110111100000010;
		b = 32'b11101011110001001101111110000011;
		correct = 32'b01010101011111111111110010011011;
		#400 //-3.695569e-14 * -4.7600993e+26 = 17591275000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010101011101101111011110000010;
		b = 32'b01001101010011000011010101110100;
		correct = 32'b11100011010001010000000011001101;
		#400 //-16971431000000.0 * 214128450.0 = -3.6340663e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110000100001111110110011010101;
		b = 32'b00000111000000011010110111010011;
		correct = 32'b00111000000010011011010101000101;
		#400 //3.365343e+29 * 9.755964e-35 = 3.2832166e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001010011001001100110011011110;
		b = 32'b10110011110110001000110010111100;
		correct = 32'b10111110110000011000101010100011;
		#400 //3748663.5 * -1.0083883e-07 = -0.37801084
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101110101100100010011101000010;
		b = 32'b00111100010111011110000001011001;
		correct = 32'b00101011100110100110100000000100;
		#400 //8.1014764e-11 * 0.013542258 = 1.0971228e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000000111111101101010110011011;
		b = 32'b01011101101011011011011101010100;
		correct = 32'b11011111001011001110110011011000;
		#400 //-7.963575 * 1.5646958e+18 = -1.2460572e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111111000101000101110111001101;
		b = 32'b10101110011111001001101100110111;
		correct = 32'b00101110000100100110011001001010;
		#400 //-0.5795563 * -5.7436025e-11 = 3.3287408e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001110000011011110010001110011;
		b = 32'b10111000110000010011000111100011;
		correct = 32'b00000111010101100010100111000010;
		#400 //-1.7489586e-30 * -9.212249e-05 = 1.6111842e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001010001110110100011000010110;
		b = 32'b11110000001111000011111101000000;
		correct = 32'b00111011000010011011010110111101;
		#400 //-9.016904e-33 * -2.3303859e+29 = 0.0021012865
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110100110011000101100100010000;
		b = 32'b01101011100000001111000100000111;
		correct = 32'b01100000110011011101100111011011;
		#400 //3.8062763e-07 * 3.1176145e+26 = 1.1866502e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010101111000000000110100100010;
		b = 32'b10111111101111011011010110100011;
		correct = 32'b11010110001001100000100010101010;
		#400 //30793376000000.0 * -1.4821056 = -45639036000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010101111111111111100100011000;
		b = 32'b11001101111000100011010011001000;
		correct = 32'b11100100011000100010111010101110;
		#400 //35180664000000.0 * -474388740.0 = -1.6689311e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111000110101010110100010110011;
		b = 32'b10100101010111000100001111000000;
		correct = 32'b01011110101101111001111001110100;
		#400 //-3.4627587e+34 * -1.9104913e-16 = 6.61557e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001011001011100100010101100011;
		b = 32'b01110110100011101011011100100001;
		correct = 32'b01000010010000100100111001001110;
		#400 //3.3563382e-32 * 1.4473056e+33 = 48.57647
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111111110010011000010100110001;
		b = 32'b11111100001110111100000011100001;
		correct = 32'b01111111110010011000010100110001;
		#400 //nan * -3.8994862e+36 = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110010000111001100110100000000;
		b = 32'b00101011001011101001011010001010;
		correct = 32'b11011101110101011101111100010101;
		#400 //-3.1057594e+30 * 6.2026133e-13 = -1.9263824e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111011101000000001010100100100;
		b = 32'b00001111101011000001100000110011;
		correct = 32'b11001011110101110011101010101100;
		#400 //-1.6623926e+36 * 1.696983e-29 = -28210520.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011010001100111111110100101000;
		b = 32'b00110000010110101111110100000110;
		correct = 32'b10001011000110011111011101111001;
		#400 //-3.722083e-23 * 7.9667506e-10 = -2.9652906e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111101110010000001011100010010;
		b = 32'b10110111110111000100000100101001;
		correct = 32'b01110110001011000010011011000001;
		#400 //-3.3245673e+37 * -2.6256386e-05 = 8.729112e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000101100101110010100111101110;
		b = 32'b11101000011011001001001110001101;
		correct = 32'b01101110100010111011000111001000;
		#400 //-4837.241 * -4.4688013e+24 = 2.161667e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100001001100110011111011110101;
		b = 32'b01001100000111001011111101111111;
		correct = 32'b10101101110110111000000011100100;
		#400 //-6.073088e-19 * 41090556.0 = -2.4954656e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011101011111001001000011101100;
		b = 32'b01010011111100101100011011101010;
		correct = 32'b11110001111011111000010100111110;
		#400 //-1.1374566e+18 * 2085438600000.0 = -2.3720959e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000011110000000000011000010010;
		b = 32'b10111100111111100100100110101010;
		correct = 32'b10000001001111101011110101000111;
		#400 //1.1286139e-36 * -0.031040985 = -3.5033288e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000001101111001000101011011011;
		b = 32'b01000010001000111100101000101101;
		correct = 32'b01000100011100010100001010100000;
		#400 //23.5678 * 40.947437 = 965.041
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000101110100110101001111011101;
		b = 32'b10111100101101011011111111000100;
		correct = 32'b10000011000101100000100010011001;
		#400 //1.9873151e-35 * -0.022186168 = -4.409091e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011101110111110111001011010011;
		b = 32'b10111010011001000100011100000111;
		correct = 32'b01011000110001110100000001000011;
		#400 //-2.0126455e+18 * -0.00087080937 = 1752630500000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011101100111001011111101010110;
		b = 32'b01110101011011101100001010001010;
		correct = 32'b11010011100100100011000011111111;
		#400 //-4.1490693e-21 * 3.0266415e+32 = -1255774500000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110110001110100101101011100010;
		b = 32'b00001111000111110011100100010001;
		correct = 32'b01000101111001111100111111111010;
		#400 //9.449322e+32 * 7.850296e-30 = 7417.997
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001100101111001111001100101001;
		b = 32'b00010100011111000110101001101100;
		correct = 32'b00100001101110100100110111101001;
		#400 //99064136.0 * 1.2743737e-26 = 1.2624473e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000000110010011111010110010100;
		b = 32'b11001101101110001111100100111100;
		correct = 32'b00001111000100011110110100100010;
		#400 //-1.8547032e-38 * -387917700.0 = 7.194722e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001010100110110000000110101001;
		b = 32'b00000001101011111111000011010010;
		correct = 32'b00001100110101010000111111100110;
		#400 //5079252.5 * 6.463041e-38 = 3.2827415e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101010101100110110000011110010;
		b = 32'b00110101000001000101000011010000;
		correct = 32'b01100000001110010110110100111010;
		#400 //1.0842777e+26 * 4.929143e-07 = 5.3445598e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011011011111100110100110010111;
		b = 32'b11010000100011100010100010111010;
		correct = 32'b01101100100011010100011100001011;
		#400 //-7.161074e+16 * -19080270000.0 = 1.3663523e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010101110100101110010110010101;
		b = 32'b01111101100100101000010011101101;
		correct = 32'b11010011111100010110100011100001;
		#400 //-8.518054e-26 * 2.4344685e+37 = -2073693400000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111000011111011010111011100001;
		b = 32'b01111000001001001011111100100000;
		correct = 32'b01110001001000110100000101101101;
		#400 //6.048277e-05 * 1.3365831e+34 = 8.084024e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011111100111101000100111001100;
		b = 32'b10110110110101101101010101011011;
		correct = 32'b01010111000001010000101101010010;
		#400 //-2.2847772e+19 * -6.402535e-06 = 146283670000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101011001001001010100101101100;
		b = 32'b00111110000101101010110000100111;
		correct = 32'b01101001110000011101010000000000;
		#400 //1.990639e+26 * 0.14714108 = 2.9290478e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101000110111111000001100110011;
		b = 32'b10001100010001000101111010110100;
		correct = 32'b10110101101010110111001100100010;
		#400 //8.4440634e+24 * -1.512779e-31 = -1.2774001e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010110101001000011110000011000;
		b = 32'b11111111111111001011001100111001;
		correct = 32'b11111111111111001011001100111001;
		#400 //-2.6533553e-25 * nan = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001100111000001110111011100111;
		b = 32'b01111101110001111101111011011011;
		correct = 32'b01001011001011111001110110000101;
		#400 //3.4656449e-31 * 3.3209188e+37 = 11509125.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000111101111100000011110010111;
		b = 32'b11000010110000001111000010111101;
		correct = 32'b10001011000011110011100001100101;
		#400 //2.8592484e-34 * -96.47019 = -2.7583225e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011100111101110100001111011011;
		b = 32'b00110010110110011111101110110000;
		correct = 32'b10010000010100101000101110011110;
		#400 //-1.6362629e-21 * 2.5376579e-08 = -4.1522755e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100111100011011000100100010001;
		b = 32'b00011100010000100011101001011011;
		correct = 32'b01000100010101101100010001000100;
		#400 //1.3367642e+24 * 6.426464e-22 = 859.06665
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010011010000101101011111010101;
		b = 32'b01101000011001101101001101111101;
		correct = 32'b11111100001011111010111011100000;
		#400 //-836844700000.0 * 4.3601822e+24 = -3.6487953e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010010010110010100111001101001;
		b = 32'b10100010101011110100101100010000;
		correct = 32'b00110101100101001100110001010001;
		#400 //-233330850000.0 * -4.751332e-18 = 1.1086323e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000000011111000001001110001111;
		b = 32'b01000100101011001011100101011101;
		correct = 32'b00000101101001110110110111110111;
		#400 //1.1394618e-38 * 1381.7926 = 1.5744999e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111000011101001100001001110011;
		b = 32'b10010000110101101110010110000010;
		correct = 32'b10001001110011010111010111111010;
		#400 //5.835523e-05 * -8.476173e-29 = -4.94629e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111001101011001000100100010110;
		b = 32'b01110011111110010001011101011111;
		correct = 32'b11101110001001111110000100010111;
		#400 //-0.00032908533 * 3.947009e+31 = -1.2989028e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110011110100011100100001001110;
		b = 32'b10101001010010001011010110000100;
		correct = 32'b10011101101001000111100100111100;
		#400 //9.768756e-08 * -4.456636e-14 = -4.353579e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001010010011001111100110110000;
		b = 32'b11001011100000011011101100000011;
		correct = 32'b00010110010011111011111100011101;
		#400 //-9.869204e-33 * -17004038.0 = 1.6781632e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110001010001111111001010001010;
		b = 32'b00101010000111000111011110100111;
		correct = 32'b10011011111101000110101010000001;
		#400 //-2.9096179e-09 * 1.3897096e-13 = -4.043524e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000110010010011110100001100000;
		b = 32'b01101111011001010110110001011101;
		correct = 32'b01110110001101001111001001010101;
		#400 //12922.094 * 7.100307e+28 = 9.175083e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100110011011000000010000011101;
		b = 32'b00100001110010011111111101001001;
		correct = 32'b11001000101110100011101010010110;
		#400 //-2.786386e+23 * 1.3687863e-18 = -381396.7
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111000100010110100101010111110;
		b = 32'b11011011000011101111011001000101;
		correct = 32'b11010100000110111001001011101010;
		#400 //6.641958e-05 * -4.0240223e+16 = -2672739000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010011000100001110111010001011;
		b = 32'b11011011101001111001110100001110;
		correct = 32'b10101111001111011100100100001110;
		#400 //1.8292966e-27 * -9.435801e+16 = -1.7260879e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011101000010000101101000000001;
		b = 32'b11001011001011000110100010111111;
		correct = 32'b11101000101101111010100010000110;
		#400 //6.140729e+17 * -11299007.0 = -6.938414e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101110001111001100000110111101;
		b = 32'b00001010000011110110001111001100;
		correct = 32'b00111000110100110111001110011100;
		#400 //1.4604349e+28 * 6.903969e-33 = 0.00010082798
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000000011101110111111011110000;
		b = 32'b01010001011110110001011100011100;
		correct = 32'b00010010011010100110100001111110;
		#400 //1.097396e-38 * 67401530000.0 = 7.3966177e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100110111010100111000010001101;
		b = 32'b01010101010110100101000101111101;
		correct = 32'b10111100110001111110111001111000;
		#400 //-1.6267519e-15 * 15002720000000.0 = -0.024405703
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110011011100100011011000000110;
		b = 32'b00011011011101001100100111100000;
		correct = 32'b01001111011001111001101001111110;
		#400 //1.9189935e+31 * 2.0248436e-22 = 3885661700.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101011101100110010111101001011;
		b = 32'b10111011011101101001001011011000;
		correct = 32'b00100111101011001001011000111010;
		#400 //-1.2731841e-12 * -0.0037624147 = 4.7902466e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001001110001100111011000100100;
		b = 32'b00110111010011111000001001110010;
		correct = 32'b00000001101000001101111010100111;
		#400 //4.7777865e-33 * 1.2368533e-05 = 5.909421e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101110101110011111010010011110;
		b = 32'b00011111001001011110111000001010;
		correct = 32'b11001110011100010000111100100101;
		#400 //-2.8775225e+28 * 3.513701e-20 = -1011075400.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100010111111011100101100011000;
		b = 32'b01010000000000100000110000001010;
		correct = 32'b10110011100000001110110100010010;
		#400 //-6.879082e-18 * 8727308000.0 = -6.003587e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011001011101001111101010110100;
		b = 32'b11100100000010011010000000100101;
		correct = 32'b10111110000000111011001101101010;
		#400 //1.26651334e-23 * -1.0154974e+22 = -0.1286141
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101101000100110100110011011111;
		b = 32'b10101111101101110011111100101101;
		correct = 32'b10011101010100101110000010011010;
		#400 //8.373051e-12 * -3.3332395e-10 = -2.7909385e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000000100100011010110111110110;
		b = 32'b10101101001100110001101111111010;
		correct = 32'b10101110010010111101100100011101;
		#400 //4.5524855 * -1.0181184e-11 = -4.634969e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010101010101000000111100010011;
		b = 32'b10011110110111011000100011010101;
		correct = 32'b00110100101101111000001001011100;
		#400 //-14572576000000.0 * -2.3455878e-20 = 3.4181255e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001001001000010001101011111111;
		b = 32'b00100010000001111010000101011110;
		correct = 32'b10101011101010101011010110010011;
		#400 //-659887.94 * 1.8381339e-18 = -1.2129623e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000100100100011101011110001100;
		b = 32'b01000110110010100111100001001011;
		correct = 32'b10001011111001101011000100111000;
		#400 //-3.4287285e-36 * 25916.146 = -8.8859427e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101111010110010110000111001000;
		b = 32'b00000011000010001011110110110010;
		correct = 32'b00110010111010000011101000001101;
		#400 //6.7276457e+28 * 4.0184567e-37 = 2.7034753e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000011111101011111101001100011;
		b = 32'b01010000110100011011000110000000;
		correct = 32'b10010101010010010111101111111000;
		#400 //-1.4457292e-36 * 28144566000.0 = -4.068942e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101100111011000111111111010010;
		b = 32'b01110100111011111000011111110010;
		correct = 32'b11100010010111010100100011101100;
		#400 //-6.7217143e-12 * 1.5182083e+32 = -1.02049625e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000101010100001101000010101;
		b = 32'b11100110001110111011101001100100;
		correct = 32'b01010111011110010111100111001101;
		#400 //-1.2376541e-09 * -2.216302e+23 = 274301530000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001011111010001000011110000100;
		b = 32'b01100100000111001010110001010100;
		correct = 32'b00110000100011100100111100011100;
		#400 //8.956705e-32 * 1.1560439e+22 = 1.0354344e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100111001110000011111001100111;
		b = 32'b00110101000101011101011001110110;
		correct = 32'b01011100110101111010110101010110;
		#400 //8.7006655e+23 * 5.581891e-07 = 4.8566164e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000000000100101011110000001010;
		b = 32'b00001101011010000110110010111111;
		correct = 32'b10001110000001010011100010111110;
		#400 //-2.292727 * 7.162142e-31 = -1.6420836e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010000111001100110001011010111;
		b = 32'b11111101111001010011100110100100;
		correct = 32'b11001111010011100100101001001010;
		#400 //9.087129e-29 * -3.8086562e+37 = -3460975000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001010100110110011111111111101;
		b = 32'b01000110111001010001111110101111;
		correct = 32'b01010010000010101111001101110100;
		#400 //5087230.5 * 29327.842 = 149197490000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101011000111000110101010011001;
		b = 32'b01000100000011101000101010111011;
		correct = 32'b01101111101011100010111111001001;
		#400 //1.8909582e+26 * 570.16766 = 1.0781632e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111011001110111111100001101101;
		b = 32'b11001111010011100000010010111110;
		correct = 32'b11001011000101110100010101100011;
		#400 //0.002868201 * -3456417300.0 = -9913699.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100100101011101111110111111100;
		b = 32'b11011011000100000011010111001100;
		correct = 32'b01000000010001010010011101001000;
		#400 //-7.589074e-17 * -4.0591547e+16 = 3.0805225
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101001011101101000110011101011;
		b = 32'b01100101010100011101010100100010;
		correct = 32'b01001111010010100001011001010000;
		#400 //5.47452e-14 * 6.1931638e+22 = 3390460000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111111110000000001001110000;
		b = 32'b01101111101111000111010010111111;
		correct = 32'b11101000001101101001001011100100;
		#400 //-2.9565039e-05 * 1.1664864e+29 = -3.4487214e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001100111001011001111100110001;
		b = 32'b11001110010111111000011001010100;
		correct = 32'b10011011110010000111111000101000;
		#400 //3.5378846e-31 * -937530600.0 = -3.316875e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100001111100000011001000011;
		b = 32'b11110101000000111011000101001110;
		correct = 32'b11111001110000111000000110100001;
		#400 //760.09784 * -1.669402e+32 = -1.2689088e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110101111101011010000111111110;
		b = 32'b00101010000010101001000010011110;
		correct = 32'b00100000100001001111010000010110;
		#400 //1.8301068e-06 * 1.2307036e-13 = 2.2523192e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100110101111010100101100000000;
		b = 32'b10100001100100110011101110001100;
		correct = 32'b10001000110110011011110000110010;
		#400 //1.3134838e-15 * -9.976869e-19 = -1.3104457e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111010011001010111101101010001;
		b = 32'b11001111011001111001001100111101;
		correct = 32'b11001010010011111001011001000011;
		#400 //0.00087540323 * -3885186300.0 = -3401104.8
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000101001011100011000010110100;
		b = 32'b11100011110111010000100000100011;
		correct = 32'b10101001100101100110010110010101;
		#400 //8.190386e-36 * -8.1546335e+21 = -6.67896e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101110111011000110010111000001;
		b = 32'b01001010000110101001101011110101;
		correct = 32'b00111001100011101100010001001110;
		#400 //1.07501126e-10 * 2533053.2 = 0.0002723061
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100011000111100001010011011110;
		b = 32'b00001011011110010110100000101101;
		correct = 32'b00101111000110100000001010100000;
		#400 //2.9160892e+21 * 4.803403e-32 = 1.4007151e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101111010110100100100001110000;
		b = 32'b10011111001000010110010010001010;
		correct = 32'b10001111000010011001110101001000;
		#400 //1.985272e-10 * -3.417624e-20 = -6.784913e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000100101001101010100110101111;
		b = 32'b01000000101111111111110001000011;
		correct = 32'b00000101111110011111100110101000;
		#400 //3.9182242e-36 * 5.9995437 = 2.3507557e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110100101111111110111111010010;
		b = 32'b10111001000100100100001000000110;
		correct = 32'b11101110010110110101000010001100;
		#400 //1.216544e+32 * -0.0001394824 = -1.6968648e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100010111000010000100110010101;
		b = 32'b10011110011111010011011110100111;
		correct = 32'b10000001110111101001011101100100;
		#400 //6.0996518e-18 * -1.3405217e-20 = -8.1767155e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010101100101000101101010000010;
		b = 32'b00101101100000010101000101010101;
		correct = 32'b11000011100101011110000101111011;
		#400 //-20389556000000.0 * 1.470172e-11 = -299.76157
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101001110111001001111101001100;
		b = 32'b00110010011011111100110111001101;
		correct = 32'b01011100110011101010101000010100;
		#400 //3.3339492e+25 * 1.3958425e-08 = 4.653668e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000101001010010101001101001110;
		b = 32'b10001101000101001001100111001010;
		correct = 32'b00010010110001001001001111000011;
		#400 //-2709.2065 * -4.579114e-31 = 1.2405765e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000110001110111011101010100010;
		b = 32'b10011111001101011001110001110100;
		correct = 32'b10100110000001010010110110101111;
		#400 //12014.658 * -3.8457656e-20 = -4.6205557e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000110111000011011001011101011;
		b = 32'b00011111000100011100000001001100;
		correct = 32'b00100110100000000111111111100000;
		#400 //28889.459 * 3.086401e-20 = 8.916445e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011011100000111111101001001010;
		b = 32'b00101111001011010000010110100111;
		correct = 32'b00001011001100100110011000011100;
		#400 //2.1833878e-22 * 1.5736266e-10 = 3.4358372e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010101001110010010011001100111;
		b = 32'b10001011001011000111001100001001;
		correct = 32'b00100000111110010111001000000000;
		#400 //-12723412000000.0 * -3.3212538e-32 = 4.225768e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111000011111001010000111110110;
		b = 32'b00111001010100011100111101010000;
		correct = 32'b10110010010011110000110011010000;
		#400 //-6.023232e-05 * 0.00020009023 = -1.2051899e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011100111011110001010001010101;
		b = 32'b10111110110001000111110011100000;
		correct = 32'b10011100001101111000000000110000;
		#400 //1.5820949e-21 * -0.38376522 = -6.07153e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111001101010000000100000010;
		b = 32'b11011100011000000000010001010011;
		correct = 32'b11100100000111100110001111110000;
		#400 //46337.008 * -2.522206e+17 = -1.1687147e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110011010000110000010011100000;
		b = 32'b01010001111100001010001001011010;
		correct = 32'b11000101101101110101000001000000;
		#400 //-4.540641e-08 * 129189495000.0 = -5866.0312
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000011100011111010110101011101;
		b = 32'b10100100110010111110011111100011;
		correct = 32'b10101000111001001110000100111011;
		#400 //287.3544 * -8.843005e-17 = -2.5410763e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101011011011101010001000001111;
		b = 32'b10011001011111010001100001110010;
		correct = 32'b10000101011010111110110011110010;
		#400 //8.4779487e-13 * -1.308473e-23 = -1.1093167e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010011111000001110100110001011;
		b = 32'b10111101100010001001010111001111;
		correct = 32'b11010001111011111111111101011111;
		#400 //1931981800000.0 * -0.06669199 = -128847700000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100000000100010100110110010110;
		b = 32'b11010100100001000001101101111110;
		correct = 32'b10110101000101011111011100111000;
		#400 //1.2307649e-19 * -4539175400000.0 = -5.5866576e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011101101010010101001000111100;
		b = 32'b10011101100100101111011100001100;
		correct = 32'b00111011110000100110100010011001;
		#400 //-1.52511e+18 * -3.890132e-21 = 0.005932879
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111110011110110000010010011010;
		b = 32'b00001101111100101110011110110110;
		correct = 32'b01001100111011100010110110001101;
		#400 //8.341503e+37 * 1.4970184e-30 = 124873830.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011101100011101101101001111101;
		b = 32'b01010010100110110101100101001101;
		correct = 32'b01110000101011010110000000111101;
		#400 //1.2867097e+18 * 333609070000.0 = 4.29258e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101100101110100101111000001001;
		b = 32'b10111010001010010000010000001100;
		correct = 32'b10100111011101100001011000001100;
		#400 //5.296878e-12 * -0.00064474414 = -3.415131e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100111111010010111000011010100;
		b = 32'b11001110010010111100111000111011;
		correct = 32'b11110110101110011101100010000111;
		#400 //2.2047854e+24 * -854822600.0 = -1.8847004e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011000011011000001000001000010;
		b = 32'b10010101011111000001110111100001;
		correct = 32'b00101110011010000111101110001110;
		#400 //-1038218300000000.0 * -5.0914565e-26 = 5.286043e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101001010001000110101001100100;
		b = 32'b10011010011101011100101110010010;
		correct = 32'b01000100001111001001011000000010;
		#400 //-1.4840742e+25 * -5.0829255e-23 = 754.3439
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010000000000001000101101110101;
		b = 32'b11111101010111100010010001111010;
		correct = 32'b11001101110111110001011010000001;
		#400 //2.5350983e-29 * -1.8454876e+37 = -467849250.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011100101111001100101100110100;
		b = 32'b10101110111000111100111100101010;
		correct = 32'b10001100001010000000000011110110;
		#400 //1.2493323e-21 * -1.03595646e-10 = -1.2942538e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100010101101011001100000101100;
		b = 32'b11000110000010001010101000000000;
		correct = 32'b11101001010000011110001011011101;
		#400 //1.6749129e+21 * -8746.5 = -1.4649626e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110001110000000000100011010100;
		b = 32'b10100110101001100101010010110001;
		correct = 32'b10011000111110011000101010000010;
		#400 //5.588939e-09 * -1.154152e-15 = -6.450485e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001111100110101010001111100011;
		b = 32'b10110100010001101010000110011110;
		correct = 32'b01000100011011111111100011000100;
		#400 //-5188863500.0 * -1.8498983e-07 = 959.88696
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010011100111110111000001010101;
		b = 32'b10000010000110011000010100110011;
		correct = 32'b10010110001111110011101000110000;
		#400 //1369568800000.0 * -1.1278891e-37 = -1.5447218e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101101101000011001010010111001;
		b = 32'b11001010100110110000110100010010;
		correct = 32'b10111000110000111011101010011000;
		#400 //1.8369627e-11 * -5080713.0 = -9.3330804e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110001010000010111000011110011;
		b = 32'b01110000100000000010000111011100;
		correct = 32'b11100010010000011010010000011111;
		#400 //-2.81494e-09 * 3.172401e+29 = -8.9301194e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000100111100110001011001100110;
		b = 32'b10110011111111011111010111111101;
		correct = 32'b00111001011100010010011010110111;
		#400 //-1944.7 * -1.18259756e-07 = 0.00022997973
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010010100010011111100101111010;
		b = 32'b01000110111100000100010111100101;
		correct = 32'b01011010000000010111111110001110;
		#400 //296298020000.0 * 30754.947 = 9112630000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101011111000000011101001001111;
		b = 32'b11001111110001000111100100100000;
		correct = 32'b01111100001011000001011010111100;
		#400 //-5.4214948e+26 * -6592545000.0 = 3.5741447e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101001110010100110000000001101;
		b = 32'b10101111111100001111011111011001;
		correct = 32'b10011010001111100111110111111010;
		#400 //8.987264e-14 * -4.3831852e-10 = -3.9392842e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111010011001110010111110010100;
		b = 32'b00110100100011110111000010101100;
		correct = 32'b11101111100000011000100101010100;
		#400 //-3.000964e+35 * 2.6717805e-07 = -8.017917e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011011100000100001100111100001;
		b = 32'b11011001010101111001000011111110;
		correct = 32'b11110101010110110001101011010111;
		#400 //7.32404e+16 * -3792283800000000.0 = -2.7774839e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011100001110101100001100111001;
		b = 32'b00111111110010000111101001000001;
		correct = 32'b01011100100100100100000110110101;
		#400 //2.1027598e+17 * 1.5662309 = 3.2934074e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011010001111101110000110001011;
		b = 32'b01100001001100100010100001011110;
		correct = 32'b01111100000001001101011011101100;
		#400 //1.3432058e+16 * 2.0540183e+20 = 2.7589693e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010011101000101000001000000101;
		b = 32'b11011011110011110100110000011011;
		correct = 32'b10110000000000111001011101110010;
		#400 //4.102276e-27 * -1.16698e+17 = -4.787274e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101001011001110111101101101100;
		b = 32'b10111100111110111111001111011101;
		correct = 32'b10100110111000111101001010000101;
		#400 //5.1399355e-14 * -0.030755932 = -1.5808351e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100101001110111010101101001001;
		b = 32'b11000000100011001011101010000001;
		correct = 32'b11100110010011100101010011001010;
		#400 //5.5390137e+22 * -4.3977666 = -2.435929e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010011001010010100110001011011;
		b = 32'b11111100000100010000001001110111;
		correct = 32'b11001111101111111100101111000010;
		#400 //2.1368445e-27 * -3.011732e+36 = -6435603500.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110011111110000010111001010001;
		b = 32'b00011000001100000011000000000010;
		correct = 32'b11001100101010101100111001100010;
		#400 //-3.9325837e+31 * 2.2771705e-24 = -89551630.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000011010100100110100001111;
		b = 32'b00111110110100011110000110010110;
		correct = 32'b10101111110000000001011101100000;
		#400 //-8.523821e-10 * 0.4099242 = -3.4941205e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011111011000001011100101110111;
		b = 32'b01000110001011100100011110010110;
		correct = 32'b00100110000110001111110011100110;
		#400 //4.7587258e-20 * 11153.896 = 5.3078335e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000111110001101110010110101100;
		b = 32'b10111110111011101101010001110001;
		correct = 32'b10000111001110011000111010010100;
		#400 //2.9926718e-34 * -0.46646455 = -1.3959753e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111100101001110010011101010010;
		b = 32'b11101000101101110110100111001111;
		correct = 32'b11100101111011111000010001100100;
		#400 //0.020404492 * -6.929159e+24 = -1.4138597e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110101001001110000110111001101;
		b = 32'b11111100100010010110001100101101;
		correct = 32'b01110010001100110100111000110101;
		#400 //-6.223243e-07 * -5.7068495e+36 = 3.5515112e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100010011111101111100000100010;
		b = 32'b10110101001001001000011001111100;
		correct = 32'b01011000001000111101110011100111;
		#400 //-1.1758382e+21 * -6.129046e-07 = 720676650000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011101010100000100110000111011;
		b = 32'b11001011011100010010111100001100;
		correct = 32'b00101001010001000011111000001011;
		#400 //-2.7567981e-21 * -15806220.0 = 4.3574556e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001100001101000010101011110110;
		b = 32'b11011010001010011100000011110001;
		correct = 32'b10100110111011101111000001001100;
		#400 //1.3879624e-31 * -1.1945353e+16 = -1.65797e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000110110101110001001010010111;
		b = 32'b01101000011111111001101111100111;
		correct = 32'b01101111110101101011111001111111;
		#400 //27529.295 * 4.8283174e+24 = 1.3292018e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100111111100011110001101111111;
		b = 32'b01011100011010001110010010100000;
		correct = 32'b01000100110111000000111000110001;
		#400 //6.713759e-15 * 2.6221428e+17 = 1760.4435
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010001010011100110010100110101;
		b = 32'b10001010100100010000101011011100;
		correct = 32'b00011100011010011110000000101001;
		#400 //-55403827000.0 * -1.3967077e-32 = 7.7382953e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110000010100110101011100010111;
		b = 32'b11000000110110011011000110111001;
		correct = 32'b01110001101100111011011110001010;
		#400 //-2.6162649e+29 * -6.8029447 = 1.7798305e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101000001000101010111010111010;
		b = 32'b01010001011010100000100100101000;
		correct = 32'b00111010000101001011100110001000;
		#400 //9.030694e-15 * 62823498000.0 = 0.0005673398
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101111111100111001010110111001;
		b = 32'b11101100011010110011110001011100;
		correct = 32'b01011100110111111101001111011111;
		#400 //-4.4307827e-10 * -1.1375304e+27 = 5.04015e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100010110011001010110011000000;
		b = 32'b10101111010100111111001100010100;
		correct = 32'b00010010101010010111010010111010;
		#400 //-5.5477217e-18 * -1.9276697e-10 = 1.0694175e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100001100001011011100110100101;
		b = 32'b10100000111010110101100110010011;
		correct = 32'b11000010111101011110000001101010;
		#400 //3.0834926e+20 * -3.9869824e-19 = -122.93831
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000011100010001111010110010001;
		b = 32'b10100100010101001011010101001011;
		correct = 32'b00101000011000111001100010110100;
		#400 //-273.9185 * -4.6123733e-17 = 1.26341435e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101111100110101101010011011100;
		b = 32'b01001100010000010100000011100111;
		correct = 32'b11111100011010011100001101110110;
		#400 //-9.583605e+28 * 50660252.0 = -4.8550783e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010000111011001000011110101010;
		b = 32'b01011010110100010100011000111010;
		correct = 32'b00101100010000010101101110100100;
		#400 //9.329461e-29 * 2.9452743e+16 = 2.747782e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111011010000001101111101001100;
		b = 32'b00011001011010110111101001010101;
		correct = 32'b01010101001100010110100100100101;
		#400 //1.00145e+36 * 1.217392e-23 = 12191572000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110110110011010110110010101000;
		b = 32'b10111010101011001110100101000010;
		correct = 32'b01110010000010101100000000101110;
		#400 //-2.0832513e+33 * -0.0013192075 = 2.7482408e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110111110100010100110000000110;
		b = 32'b10111011101001000010101101001100;
		correct = 32'b10110100000001100011100000011010;
		#400 //2.4950143e-05 * -0.005010044 = -1.2500132e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001110100001101011000100101000;
		b = 32'b11000101000100110010101110010001;
		correct = 32'b10010100000110101101110101001100;
		#400 //3.3204146e-30 * -2354.723 = -7.818656e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011101101101000001011111100000;
		b = 32'b10110101111110001111101001111111;
		correct = 32'b10010100001011110010011101011010;
		#400 //4.767029e-21 * -1.8550344e-06 = -8.843003e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011101001000111001110101010111;
		b = 32'b10110001111001111110101011011111;
		correct = 32'b01001111100101000011100100010110;
		#400 //-7.368547e+17 * -6.7496866e-09 = 4973538300.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101100000111101001101101010000;
		b = 32'b11100100101011011101000111111100;
		correct = 32'b11010001010101110110001000011100;
		#400 //2.2539366e-12 * -2.5651342e+22 = -57816500000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101111010111111010111011110010;
		b = 32'b10110101100000101110111101010111;
		correct = 32'b00100101011001001100111111101110;
		#400 //-2.0343885e-10 * -9.755412e-07 = 1.9846297e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000000101101001100111010110110;
		b = 32'b10011111001110101110111110110111;
		correct = 32'b10100000100001000000011101111110;
		#400 //5.6502333 * -3.958532e-20 = -2.2366628e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001110000010100111111101100101;
		b = 32'b01000011010001110111111100111011;
		correct = 32'b00010001110101111101101110111001;
		#400 //1.7071152e-30 * 199.497 = 3.4056433e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000101100101100111111011110111;
		b = 32'b11010010011100000011011010101101;
		correct = 32'b00011000100011010011011100101100;
		#400 //-1.4152572e-35 * -257927360000.0 = 3.6503355e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111100011011101101111011101000;
		b = 32'b10001000110001000001100001010111;
		correct = 32'b11000101101101101111100101100000;
		#400 //4.961151e+36 * -1.1802043e-33 = -5855.172
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001111100000101110111011000101;
		b = 32'b10010111001111110100111100000010;
		correct = 32'b00100111010000111011000100011011;
		#400 //-4393372000.0 * -6.181515e-25 = 2.7157695e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010100001110010001100101011101;
		b = 32'b00010011001101111001011011011111;
		correct = 32'b10101000000001001011111000111000;
		#400 //-3179978000000.0 * 2.3172232e-27 = -7.368719e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101110001110111100101111110100;
		b = 32'b10101101010010100111001111001101;
		correct = 32'b01011100000101001000001111100010;
		#400 //-1.4530065e+28 * -1.15080835e-11 = 1.6721321e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100110000101110111011011100101;
		b = 32'b11100111101110110100110100100000;
		correct = 32'b01001110010111011010001011110110;
		#400 //-5.254978e-16 * -1.7690105e+24 = 929611140.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110100000100000011100100111101;
		b = 32'b11010011101100001111101011011000;
		correct = 32'b11001000010001110110100101010111;
		#400 //1.3431868e-07 * -1520245400000.0 = -204197.36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100010110000100011010011010100;
		b = 32'b01010010001100110110010001100001;
		correct = 32'b11110101100010000001011100010110;
		#400 //-1.7912375e+21 * 192620800000.0 = -3.450296e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011001110001001110100110110001;
		b = 32'b00100111100100000010101000000010;
		correct = 32'b11000001110111011100011110000111;
		#400 //-6928255000000000.0 * 4.0013574e-15 = -27.722425
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000001011100011100000101011010;
		b = 32'b00110011101111011011110111001001;
		correct = 32'b00110101101100110010111011111001;
		#400 //15.109705 * 8.83552e-08 = 1.335021e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010101101100001110100000100010;
		b = 32'b11001101111101010111011110110111;
		correct = 32'b00100100001010011010000011100011;
		#400 //-7.1452075e-26 * -514782940.0 = 3.678231e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011101010010010111100100001011;
		b = 32'b01111101101100001110101101100011;
		correct = 32'b01011011100010110011110001111000;
		#400 //2.6664706e-21 * 2.939579e+37 = 7.838302e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000011000111100110111010011000;
		b = 32'b00111100111101110000000111010100;
		correct = 32'b11000000100110001101110111010110;
		#400 //-158.432 * 0.030152239 = -4.7770796
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100001110100001001000100111011;
		b = 32'b01011010110101000001110001000100;
		correct = 32'b10111101001011001100111101001100;
		#400 //-1.413307e-18 * 2.9851887e+16 = -0.04218988
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011011110001100101100101010001;
		b = 32'b01100111111100010010001111011000;
		correct = 32'b01000100001110101101010111011011;
		#400 //3.2814072e-22 * 2.277503e+24 = 747.3415
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010100111111101101000011001101;
		b = 32'b00110001011101000010010100111011;
		correct = 32'b10000110111100110000010000010010;
		#400 //-2.5729803e-26 * 3.5527836e-09 = -9.141242e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001111011100010000011001011010;
		b = 32'b10110011001011000011000011010001;
		correct = 32'b11000011001000100001111000111010;
		#400 //4043725300.0 * -4.009127e-08 = -162.11807
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001001100101010100001000111000;
		b = 32'b11101000000001010100010001101000;
		correct = 32'b11110010000110110110011010010011;
		#400 //1222727.0 * -2.5173465e+24 = -3.0780276e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001001110000100000010001001111;
		b = 32'b01000101001010111100000011101010;
		correct = 32'b01001111100000100010101100010101;
		#400 //1589385.9 * 2748.0571 = 4367723000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111001010010111000011101011101;
		b = 32'b01010001010011011101110010000100;
		correct = 32'b11001011001000111010101010110111;
		#400 //-0.00019410015 * 55260496000.0 = -10726071.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001100010101110001001111000111;
		b = 32'b01010100101000110111111100010100;
		correct = 32'b00100001100010010101110001011011;
		#400 //1.6568949e-31 * 5617693500000.0 = 9.307927e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001011100110001110001110110011;
		b = 32'b01100110100001001011011100111100;
		correct = 32'b01110010100111101000010110101110;
		#400 //20039526.0 * 3.1336623e+23 = 6.279711e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011000011010010010001110100111;
		b = 32'b00111001100000001010010111001110;
		correct = 32'b01010010011010100101000110100110;
		#400 //1025357340000000.0 * 0.00024537597 = 251598050000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000111011000010010100011001011;
		b = 32'b01010111111010100100000111001110;
		correct = 32'b10011111110011100000100100101010;
		#400 //-1.6939107e-34 * 515136700000000.0 = -8.7259554e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000011100010001000000011001101;
		b = 32'b01000111010011111101100111000011;
		correct = 32'b01001011010111011010100010000110;
		#400 //273.00626 * 53209.76 = 14526598.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001001000101001100000010111010;
		b = 32'b11010010011010010011111010110100;
		correct = 32'b01011100000001111000011111011001;
		#400 //-609291.6 * -250444840000.0 = 1.5259395e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010010111000011001111101001001;
		b = 32'b01010111100100100111100110010010;
		correct = 32'b00101011000000010001011111111101;
		#400 //1.4238763e-27 * 322101680000000.0 = 4.5863297e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000011011011001001000100100000;
		b = 32'b10011101001101010010101111011101;
		correct = 32'b10100001001001110110101100100100;
		#400 //236.5669 * -2.3977827e-21 = -5.67236e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110100110010010011011011001110;
		b = 32'b10010100010100001101111011001110;
		correct = 32'b10001001101001000010101110100111;
		#400 //3.7479043e-07 * -1.0545257e-26 = -3.9522614e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011000110011101011101000111;
		b = 32'b01000101010011111110001111010100;
		correct = 32'b11010000111110011101101111110111;
		#400 //-10082119.0 * 3326.2393 = -33535540000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111101100110110001100001001000;
		b = 32'b10001111101100010011111010010011;
		correct = 32'b10001101110101101100001101100101;
		#400 //0.07572991 * -1.747765e-29 = -1.3235808e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011000101001001000100001100011;
		b = 32'b01011011110001001100110101011111;
		correct = 32'b01110100111111001111100011010100;
		#400 //1447245500000000.0 * 1.1078981e+17 = 1.6034004e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000101110101010101111011011111;
		b = 32'b01010011000100110001100101111000;
		correct = 32'b11011001011101010011010101101001;
		#400 //-6827.859 * 631787500000.0 = -4313756000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101000111111100010110100100111;
		b = 32'b00110001010101010101011010001010;
		correct = 32'b00011010110100111101000101111110;
		#400 //2.8219247e-14 * 3.1044771e-09 = 8.760601e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101000010101000100010010100111;
		b = 32'b10001000100001110110100011100010;
		correct = 32'b10110001011000001000111001010111;
		#400 //4.0096324e+24 * -8.149675e-34 = -3.26772e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101010110110001001101100010011;
		b = 32'b01010110011111100010000110111100;
		correct = 32'b11000001110101110000011001101000;
		#400 //-3.8476912e-13 * 69855210000000.0 = -26.878128
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000001110100100110000110010001;
		b = 32'b01110110100101011010011111101111;
		correct = 32'b00111000111101011111100110010111;
		#400 //7.728182e-38 * 1.517692e+33 = 0.00011729
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011011111011010001001110011101;
		b = 32'b11001100100000101100110000010110;
		correct = 32'b00101000111100100100000111101011;
		#400 //-3.9221036e-22 * -68575410.0 = 2.6895985e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110111010001011001010101010;
		b = 32'b00011100100001100011101111001011;
		correct = 32'b10010011111101000000011110111101;
		#400 //-6.934938e-06 * 8.882832e-22 = -6.160189e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100001110000101010010111111000;
		b = 32'b00110101110011011100101001100100;
		correct = 32'b11011000000111000111100011001011;
		#400 //-4.4882846e+20 * 1.5332594e-06 = -688170460000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101100101111100110111111111001;
		b = 32'b00010111110110111010100110110011;
		correct = 32'b01000101001000110110100000000111;
		#400 //1.8417975e+27 * 1.4195381e-24 = 2614.5017
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010100111010000001001011110100;
		b = 32'b11001100011110101100110111111010;
		correct = 32'b11100001111000110101110100111100;
		#400 //7974003000000.0 * -65746920.0 = -5.2426614e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110001100011001111000000000100;
		b = 32'b11000110111101010001110111011001;
		correct = 32'b11111001000001101111001000100010;
		#400 //1.395778e+30 * -31374.924 = -4.3792426e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000001010100101111110011111100;
		b = 32'b11010101100111001011010101010101;
		correct = 32'b10010111100000010010011110011100;
		#400 //3.8752416e-38 * -21537829000000.0 = -8.346428e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111010101110100100000000110101;
		b = 32'b00011000010010001111111111100011;
		correct = 32'b00010011100100100011110001010101;
		#400 //0.0014209809 * 2.5978584e-24 = 3.6915073e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001000000001111011101000110010;
		b = 32'b11001110000010001100011001101101;
		correct = 32'b01010110100100010000100000111101;
		#400 //-138984.78 * -573676350.0 = 79732285000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111001101000010000001010101101;
		b = 32'b01011101000000000101110110011001;
		correct = 32'b11010111001000010111100001101001;
		#400 //-0.00030710307 * 5.7810734e+17 = -177538530000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110110110001000111101100111010;
		b = 32'b00010110100001100010111100001000;
		correct = 32'b11001101110011011111100100110010;
		#400 //-1.9925576e+33 * 2.1678548e-25 = -431957570.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011011011100101111110001111100;
		b = 32'b11000011101011111001000001110010;
		correct = 32'b01011111101001101010001110110011;
		#400 //-6.8394554e+16 * -351.12848 = 2.4015276e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010111101011000010111010000010;
		b = 32'b10000100101111011001100100101111;
		correct = 32'b10011100111111110000101010111011;
		#400 //378631500000000.0 * -4.4574363e-36 = -1.6877258e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100110000000011100100100000011;
		b = 32'b00010110001101111100100100100010;
		correct = 32'b10111100101110100101100101010010;
		#400 //-1.5322332e+23 * 1.4846089e-25 = -0.02274767
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010101101110110101000100001000;
		b = 32'b01101110010101110111111011110011;
		correct = 32'b01000100100111011010110111110001;
		#400 //7.5656543e-26 * 1.6673187e+28 = 1261.4357
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010001111000011011010101011011;
		b = 32'b10011001011101011100101011100011;
		correct = 32'b10101011110110001011010101110001;
		#400 //121176285000.0 * -1.2707176e-23 = -1.5398083e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011100010010110101011000000001;
		b = 32'b10101100000100001011110000110011;
		correct = 32'b11001000111001011110101110111000;
		#400 //2.2893593e+17 * -2.0568102e-12 = -470877.75
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011011001001100010111100010000;
		b = 32'b01001000000111000100100001010110;
		correct = 32'b01100011110010101110011101000110;
		#400 //4.677659e+16 * 160033.34 = 7.4858146e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110000011111000010100010100000;
		b = 32'b00011000000101110010001001010011;
		correct = 32'b11001001000101001101110111000110;
		#400 //-3.1215734e+29 * 1.9533622e-24 = -609756.4
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010101110011111101101001101011;
		b = 32'b01010000001001110011010001011010;
		correct = 32'b11100110100001111100000111111101;
		#400 //-28567126000000.0 * 11220904000.0 = -3.2054896e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010110000010011110100000000000;
		b = 32'b10001011011010100110010010100100;
		correct = 32'b10100001111111001000100010001110;
		#400 //37907380000000.0 * -4.5142474e-32 = -1.711233e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100000111110111110100001111100;
		b = 32'b11101101100111000000100000110111;
		correct = 32'b01001111000110011000100111000001;
		#400 //-4.26749e-19 * -6.036199e+27 = 2575942000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011001111100101000000011001101;
		b = 32'b11011111000100011001010001110101;
		correct = 32'b11111001100010011110011110010101;
		#400 //8532320300000000.0 * -1.0490138e+19 = -8.950521e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001000110001100000111000000111;
		b = 32'b10011000111100101001111111000111;
		correct = 32'b10100010001110111011010011011111;
		#400 //405616.22 * -6.2716868e-24 = -2.5438978e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110001000101111000100101000001;
		b = 32'b11000100001011110110011110110001;
		correct = 32'b00110101110011111010100001101001;
		#400 //-2.2051412e-09 * -701.6202 = 1.5471716e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101001010111001010010001110011;
		b = 32'b10100010100100101011010101111110;
		correct = 32'b01001100011111001110010001101101;
		#400 //-1.6671267e+25 * -3.976554e-18 = 66294196.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000101000001011101111001100011;
		b = 32'b01000011110000000111000101100110;
		correct = 32'b00001001010010010100010000101110;
		#400 //6.294476e-36 * 384.88593 = 2.4226553e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110011111100111111110000110111;
		b = 32'b00111010110001101111100101000010;
		correct = 32'b00101111001111011010001010100010;
		#400 //1.1361447e-07 * 0.0015180486 = 1.7247229e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000011101110011100011001011011;
		b = 32'b11110110011101010111010011001101;
		correct = 32'b01111010101100100001111110011000;
		#400 //-371.54965 * -1.2446111e+33 = 4.624348e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111000100101001111010000110101;
		b = 32'b00100100100100100111100000001010;
		correct = 32'b10011101101010100111001000111101;
		#400 //-7.102677e-05 * 6.352076e-17 = -4.5116745e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001010101111011111010001010101;
		b = 32'b01110101010100101110001100100001;
		correct = 32'b01000000100111000111101011110110;
		#400 //1.8291945e-32 * 2.6733131e+32 = 4.89001
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001111001010100001110000000000;
		b = 32'b00110001100000100111000101001100;
		correct = 32'b11000001001011010101101100000010;
		#400 //-2853961700.0 * 3.7963783e-09 = -10.834719
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011001001011101111011111110101;
		b = 32'b00111001010101100110011001000011;
		correct = 32'b00010011000100101000100100101011;
		#400 //9.045664e-24 * 0.00020446726 = 1.849542e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100001001011100110001000010110;
		b = 32'b10111010000110011111111100101001;
		correct = 32'b10011011110100011100110011011110;
		#400 //5.908331e-19 * -0.00058745086 = -3.4708542e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010101100111011000101110100001;
		b = 32'b01111110101110110000001010110111;
		correct = 32'b01010100111001100010110101010101;
		#400 //6.363209e-26 * 1.2428987e+38 = 7908824000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101100000010101100100010100001;
		b = 32'b10100111000010111111001101110011;
		correct = 32'b10010011100101111011110111010100;
		#400 //1.972235e-12 * -1.94221e-15 = -3.8304944e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001110101111110110000110101010;
		b = 32'b00110110011100110110001110011001;
		correct = 32'b11000101101101011111010000101010;
		#400 //-1605424400.0 * 3.6267795e-06 = -5822.5205
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000010111110011001001100111100;
		b = 32'b11010011011100001001110110000111;
		correct = 32'b01010110111010101001001110011011;
		#400 //-124.78757 * -1033435000000.0 = 128959840000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011011001011110001010010001000;
		b = 32'b11011000001001100001111110000000;
		correct = 32'b00110011111000110011100110110110;
		#400 //-1.4482295e-22 * -730616900000000.0 = 1.0581009e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101100110111101011110001100010;
		b = 32'b00001011101101101110001001000011;
		correct = 32'b00111001000111110001111011001010;
		#400 //2.1541692e+27 * 7.044429e-32 = 0.00015174891
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000100111000010001110010110111;
		b = 32'b01011110001110001100010011011100;
		correct = 32'b00100011101000100111100110111111;
		#400 //5.2923616e-36 * 3.328502e+18 = 1.7615637e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001000011101010111111111100100;
		b = 32'b00101111111010110100111011101100;
		correct = 32'b10111000111000011010100000010110;
		#400 //-251391.56 * 4.2802328e-10 = -0.000107601445
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101001001100000010100101110110;
		b = 32'b10011001100110101111101000101100;
		correct = 32'b10000011010101010100101000110000;
		#400 //3.9115812e-14 * -1.602427e-23 = -6.2680237e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101011001011010100110001001110;
		b = 32'b10100111110001001010111111111101;
		correct = 32'b00010011100001010010010110001110;
		#400 //-6.156784e-13 * -5.4591735e-15 = 3.361095e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011000101000010010010010010010;
		b = 32'b00100111110001100101011010011111;
		correct = 32'b01000000111110011011000110011111;
		#400 //1417427500000000.0 * 5.5049954e-15 = 7.8029323
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111110101011101000000011101000;
		b = 32'b10011011110111011100001011010001;
		correct = 32'b01011011000101110010101000010100;
		#400 //-1.159775e+38 * -3.668728e-22 = 4.2548987e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001010000110100001011000101011;
		b = 32'b11011001110100100111111011000001;
		correct = 32'b10100100011111010110010011110101;
		#400 //7.4189996e-33 * -7406139000000000.0 = -5.4946144e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100001010011001001100100001101;
		b = 32'b11001001111100010110000100101100;
		correct = 32'b00101011110000001110100110111110;
		#400 //-6.932045e-19 * -1977381.5 = 1.3707297e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010111101001011000011110000001;
		b = 32'b10101100001110001110011110111111;
		correct = 32'b00000100011011110001111001111011;
		#400 //-1.0697081e-24 * -2.6276618e-12 = 2.8108311e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101111001001010111011111110011;
		b = 32'b01001111011111011110110110110110;
		correct = 32'b11111111001001000010000100110001;
		#400 //-5.1210036e+28 * 4260214300.0 = -2.1816573e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000000001000110100011111111110;
		b = 32'b11101101010100100000110011000001;
		correct = 32'b01101110000001011111100100110001;
		#400 //-2.551269 * -4.0629544e+27 = 1.036569e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101011011001101001100101110111;
		b = 32'b00110110000000110001011101010100;
		correct = 32'b00100001111011000010101100010111;
		#400 //8.192539e-13 * 1.95341e-06 = 1.6003388e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011001101001010101101010001000;
		b = 32'b00101000101110000101100100000100;
		correct = 32'b01000010111011100010010100100010;
		#400 //5817864000000000.0 * 2.0466708e-14 = 119.072525
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011001111001111101001110011100;
		b = 32'b00101100101101111010111001110110;
		correct = 32'b10000111001001100101011001000001;
		#400 //-2.3970309e-23 * 5.220542e-12 = -1.25138e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011111010110010010101101010101;
		b = 32'b01111011011111101111001010110011;
		correct = 32'b11011011010110000100011011100001;
		#400 //-4.598738e-20 * 1.3237659e+36 = -6.0876527e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100110100111101101100001000011;
		b = 32'b10011110001100011111100110111100;
		correct = 32'b01000101010111001101110011110111;
		#400 //-3.750616e+23 * -9.421946e-21 = 3533.8103
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011111000100101110110100111110;
		b = 32'b00101011011011001111011111010001;
		correct = 32'b11001011000010000000000011110000;
		#400 //-1.0587186e+19 * 8.4187957e-13 = -8913136.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111100100011010110111111001100;
		b = 32'b10111101000111010100110000010110;
		correct = 32'b01111010001011011100111100110011;
		#400 //-5.875051e+36 * -0.03840264 = 2.2561746e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000110110100001101100110000110;
		b = 32'b01100001111101011101111010010110;
		correct = 32'b01101001010010001001010111000100;
		#400 //26732.762 * 5.669364e+20 = 1.5155776e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011111101000101111001001011100;
		b = 32'b11101101101010000101000110000110;
		correct = 32'b01001101110101100100010111100001;
		#400 //-6.901062e-20 * -6.5115047e+27 = 449362980.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001011010011001111010101101010;
		b = 32'b00110100110010111000111100010101;
		correct = 32'b10000000101000101111100100101001;
		#400 //-3.94736e-32 * 3.7915802e-07 = -1.4966732e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000101010010111010100010001010;
		b = 32'b00000111111010100000010011101110;
		correct = 32'b00001101101110100010101111111010;
		#400 //3258.5337 * 3.5211304e-34 = 1.1473722e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101001011000001111101001011010;
		b = 32'b10011000010000011011001101001011;
		correct = 32'b10000010001010100011101001001111;
		#400 //4.9955137e-14 * -2.5035185e-24 = -1.2506361e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010110110100011011101101011001;
		b = 32'b01000100110100100110010110111010;
		correct = 32'b11011100001011000101111100000110;
		#400 //-115301290000000.0 * 1683.179 = -1.940727e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100000000011001011000111111000;
		b = 32'b11111101111101100001110001101000;
		correct = 32'b01011110100001110100001010100001;
		#400 //-1.1917346e-19 * -4.0892198e+37 = 4.873265e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111010100110101111101001100010;
		b = 32'b10111101100001110000101111101100;
		correct = 32'b01111000101000111000001010000011;
		#400 //-4.0234604e+35 * -0.06594071 = 2.6530984e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101111010111001011010010010010;
		b = 32'b01001011101111001001011111101100;
		correct = 32'b00111011101000101001011110010101;
		#400 //2.0073035e-10 * 24719320.0 = 0.0049619176
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011111100110011101111101110000;
		b = 32'b00111111101101111101110110010111;
		correct = 32'b01011111110111010000011111010011;
		#400 //2.2175408e+19 * 1.4364499 = 3.1853861e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101110101001110001110101100001;
		b = 32'b10010101001100100000111111001101;
		correct = 32'b01000100011010000111100101111100;
		#400 //-2.5859757e+28 * -3.5959278e-26 = 929.8982
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011101110010011111110110011010;
		b = 32'b01011110111100111001010101011100;
		correct = 32'b01111101010000000011000110010010;
		#400 //1.8193699e+18 * 8.776018e+18 = 1.5966822e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011100011000000010110001100110;
		b = 32'b01010100011011000110000001110111;
		correct = 32'b01110001010011101111110101100111;
		#400 //2.5239685e+17 * 4060922800000.0 = 1.0249641e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101101111100110001101000010101;
		b = 32'b10000010100000001010000001001101;
		correct = 32'b00110000111101000100101010001000;
		#400 //-9.4045486e+27 * -1.8899918e-37 = 1.777452e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000000011101000000010011101010;
		b = 32'b11011011010011110100010001111110;
		correct = 32'b11011100010001011001000101000011;
		#400 //3.8128 * -5.834063e+16 = -2.2244115e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010111001001100001000110110111;
		b = 32'b00110101111000111111101101000001;
		correct = 32'b00001101100100111110010010110011;
		#400 //5.365985e-25 * 1.6985942e-06 = 9.114632e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001101001111001110001111001011;
		b = 32'b01011011010011100000001110011000;
		correct = 32'b01101001000110000000000111110100;
		#400 //198065330.0 * 5.7987797e+16 = 1.1485372e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110001101010010010010111110000;
		b = 32'b11101110111011011101011100110011;
		correct = 32'b11100001000111010010011001010000;
		#400 //4.9228603e-09 * -3.6804054e+28 = -1.8118122e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000110011001100011101101001100;
		b = 32'b01100001111110010010100010111110;
		correct = 32'b11101000111000000001010001010001;
		#400 //-14734.824 * 5.7452188e+20 = -8.465479e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011101101010011101111101110100;
		b = 32'b11011000110100000101001111001001;
		correct = 32'b11110111000010100011110100100111;
		#400 //1.5300787e+18 * -1832466200000000.0 = -2.8038175e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101010111011100000100001110000;
		b = 32'b10010001001110101110101011010000;
		correct = 32'b10111100101011011100110001110110;
		#400 //1.43882095e+26 * -1.474517e-28 = -0.021215659
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100100011110001001100111111100;
		b = 32'b00100000010110101110000111010011;
		correct = 32'b10000101010101001000111001101101;
		#400 //-5.3906858e-17 * 1.8540037e-19 = -9.9943516e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110000001100011000100111110001;
		b = 32'b00110101100001111000001111001011;
		correct = 32'b11100110001110111111011001001001;
		#400 //-2.1978243e+29 * 1.0096641e-06 = -2.2190642e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101000100110100010100110011101;
		b = 32'b10101011101011010110000011100011;
		correct = 32'b00010100110100001101000011101111;
		#400 //-1.7115481e-14 * -1.2319281e-12 = 2.1085043e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000111111101011010011000000111;
		b = 32'b00101101001001110011111110011100;
		correct = 32'b10110101101000000111110001011000;
		#400 //-125772.055 * 9.506975e-12 = -1.1957118e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100000000100111101000111000000;
		b = 32'b11000000111011000000011110011011;
		correct = 32'b11100001100010000100100111000001;
		#400 //4.2606023e+19 * -7.3759284 = -3.1425897e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000101111001001111100010111111;
		b = 32'b11100011011001000100000000111010;
		correct = 32'b01101001110011000010011011111100;
		#400 //-7327.0933 * -4.2104857e+21 = 3.085062e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010100100100110100010001111001;
		b = 32'b00010011101010110011111010100101;
		correct = 32'b10101000110001010000010110001101;
		#400 //-5060072000000.0 * 4.322824e-27 = -2.1873801e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011011110000110010110101110;
		b = 32'b00101001100000101101010011011110;
		correct = 32'b10110101011111011110010001011100;
		#400 //-16278958.0 * 5.810086e-14 = -9.458215e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110000010000010011100100010001;
		b = 32'b00110100000001001100011011101000;
		correct = 32'b01100100110010000110111100011100;
		#400 //2.3919838e+29 * 1.236582e-07 = 2.957884e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110110100110000111111010000;
		b = 32'b11011000100101010011100001001110;
		correct = 32'b01001111111101100000110101000000;
		#400 //-6.290131e-06 * -1312552500000000.0 = 8256127000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000000011000000010001011111010;
		b = 32'b11000101011000001001000010100000;
		correct = 32'b10000110001010001010100111010101;
		#400 //8.828755e-39 * -3593.039 = -3.172206e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100000100100001100001010101000;
		b = 32'b00111101101000010111011100011101;
		correct = 32'b11011110101101101001101110001101;
		#400 //-8.3448675e+19 * 0.07884047 = -6.579133e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101101100100000000110111010101;
		b = 32'b11000000100010100011100000101110;
		correct = 32'b00101110100110111000111000100011;
		#400 //-1.6377047e-11 * -4.319358 = 7.0738325e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000011100101100110111101000000;
		b = 32'b00011001100000101000001111101000;
		correct = 32'b10011101100110010110010000000100;
		#400 //-300.86914 * 1.3494961e-23 = -4.0602177e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100101110101110111101010001111;
		b = 32'b11100011001101010001000010011101;
		correct = 32'b01001001100110000110011110100011;
		#400 //-3.7379604e-16 * -3.3400578e+21 = 1248500.4
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100101000011100101011010001;
		b = 32'b10111010000000010110001111001010;
		correct = 32'b10111111001000111000110010001001;
		#400 //1294.338 * -0.0004935829 = -0.63886315
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010110100001011100100001000100;
		b = 32'b11011011010110101110001101001101;
		correct = 32'b10110010011001001100011010100101;
		#400 //2.1613694e-25 * -6.1611465e+16 = -1.3316513e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011101101110100110101101110010;
		b = 32'b10110001000111110110011100101110;
		correct = 32'b11001111011010000010011110111101;
		#400 //1.6791195e+18 * -2.3196196e-09 = -3894918400.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000000100100110111011100010100;
		b = 32'b01100000000000010101001011110001;
		correct = 32'b01100001000101001111110110010000;
		#400 //4.608286 * 3.7275102e+19 = 1.7177433e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001000011101111101110110010111;
		b = 32'b11000111101100011001000001101010;
		correct = 32'b01010000101010111110110000001001;
		#400 //-253814.36 * -90912.83 = 23074982000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100100011110100100110010011110;
		b = 32'b00101011000101111101000100101001;
		correct = 32'b00010000000101000110111110110010;
		#400 //5.4275006e-17 * 5.3936245e-13 = 2.92739e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011110000000100101100111101110;
		b = 32'b00101100000001011011011100010011;
		correct = 32'b10001010100010000010101111100001;
		#400 //-6.90074e-21 * 1.9002063e-12 = -1.3112829e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010001000001110111100100010001;
		b = 32'b00111000011110111011001001001000;
		correct = 32'b00001010000001010011001000001100;
		#400 //1.0686929e-28 * 6.00091e-05 = 6.41313e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011000001101111111001010000100;
		b = 32'b01010000110001000110001110001010;
		correct = 32'b01101001100011010001110100110011;
		#400 //809008900000000.0 * 26358862000.0 = 2.1324554e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000011111011001011010011101000;
		b = 32'b10000011110011001101001011010100;
		correct = 32'b10001000001111010110001100011001;
		#400 //473.41333 * -1.2038446e-36 = -5.6991607e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100101010100111010111000100001;
		b = 32'b00101100000100100001001010101000;
		correct = 32'b10010001111100011001000101111000;
		#400 //-1.836033e-16 * 2.0758204e-12 = -3.8112748e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111010000000010101010011111;
		b = 32'b10110010011000010111000000001101;
		correct = 32'b10111010001010010011100110010010;
		#400 //49194.62 * -1.3122201e-08 = -0.0006455417
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101100011011010000001111110110;
		b = 32'b00101001111111111101010011011011;
		correct = 32'b10010110111011001101110000000100;
		#400 //-3.3681924e-12 * 1.13611994e-13 = -3.8266706e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111111110000101101010010000011;
		b = 32'b01011000101111011011000000111001;
		correct = 32'b01011001000100000101110100000010;
		#400 //1.5221103 * 1668516500000000.0 = 2539666200000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100011100011101111111111000100;
		b = 32'b10111110100001100111110100101101;
		correct = 32'b01100010100101100011111110011001;
		#400 //-5.275735e+21 * -0.26267377 = 1.3857972e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110100110111110001100111011011;
		b = 32'b11011000011010010100001011000110;
		correct = 32'b01001101110010110100100010111010;
		#400 //-4.15558e-07 * -1025892000000000.0 = 426317630.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110101111110110110010111010011;
		b = 32'b10010110110001001010110100011010;
		correct = 32'b11001101010000010010001111110011;
		#400 //6.3736902e+32 * -3.177475e-25 = -202522420.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010011101111100110001110001001;
		b = 32'b01001111111000100001011011110101;
		correct = 32'b01100100001010000010010011110010;
		#400 //1635427400000.0 * 7586310700.0 = 1.2406861e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110101101111101011000111100100;
		b = 32'b11001011001111100100001110011011;
		correct = 32'b01000001100011011011101001100011;
		#400 //-1.4207876e-06 * -12469147.0 = 17.71601
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100100100010001100000010011000;
		b = 32'b01010101110001001010101110110111;
		correct = 32'b11111010110100100001111001011110;
		#400 //-2.018108e+22 * 27030224000000.0 = -5.4549913e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011010101100100010101110000000;
		b = 32'b11100010010001000000010110111011;
		correct = 32'b11111101100010000110110101001011;
		#400 //2.5075187e+16 * -9.039937e+20 = -2.266781e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011011110001010011110111001010;
		b = 32'b01010010010101000001100110100101;
		correct = 32'b01101110101000110110101011101101;
		#400 //1.1103702e+17 * 227740830000.0 = 2.528766e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011010001111100101011111010100;
		b = 32'b11001111100110111011011001100010;
		correct = 32'b01101010011001111000110110010001;
		#400 //-1.3394203e+16 * -5224842000.0 = 6.99826e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010111111110110111111101001010;
		b = 32'b11100011011000111011101011111010;
		correct = 32'b11111011110111111011100110001111;
		#400 //553048240000000.0 * -4.200884e+21 = -2.3232915e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011000111101101001001011001011;
		b = 32'b11101100101000110000011101111001;
		correct = 32'b11000110000111010000011010101010;
		#400 //6.3737733e-24 * -1.5767216e+27 = -10049.666
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010110010111111011010110110101;
		b = 32'b11001110111011101010110010010100;
		correct = 32'b11100101110100001001000110111110;
		#400 //61492880000000.0 * -2002143700.0 = -1.2311759e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010010010010011101100011010110;
		b = 32'b00110100111101011100001110111011;
		correct = 32'b00000111110000011100011011011000;
		#400 //6.369169e-28 * 4.577722e-07 = 2.9156282e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011011011110010001001100001011;
		b = 32'b01001001000000011110111110010100;
		correct = 32'b01100100111111001101011101100011;
		#400 //7.0108207e+16 * 532217.25 = 3.7312798e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011010000011011010011101101010;
		b = 32'b00110011010101010000110011100001;
		correct = 32'b11001101111010111100011011010111;
		#400 //-9968011000000000.0 * 4.960464e-08 = -494459620.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010011111101011010101110011000;
		b = 32'b11000111001000011110000111011011;
		correct = 32'b01011011100110110101100110101001;
		#400 //-2110291700000.0 * -41441.855 = 8.745441e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101101110111011101100000100001;
		b = 32'b10011000101100010111101010001001;
		correct = 32'b10000111000110011100110010011111;
		#400 //2.5220772e-11 * -4.5877157e-24 = -1.1570573e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001111000110011010100101100000;
		b = 32'b00001111000101011111100011000000;
		correct = 32'b00011110101101000000100111001000;
		#400 //2578014200.0 * 7.394175e-30 = 1.9062287e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110001110000000011101100010110;
		b = 32'b10000100000100010010100101010000;
		correct = 32'b10110110010110100000000011111010;
		#400 //1.9037617e+30 * -1.7063638e-36 = -3.24851e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000001101111111010110110000010;
		b = 32'b11100000100100000111001001110000;
		correct = 32'b01100010110110000100111010010000;
		#400 //-23.95972 * -8.326804e+19 = 1.9950789e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110110110111011100010110111001;
		b = 32'b10100011100000110101110110011101;
		correct = 32'b01011010111000111001101010001101;
		#400 //-2.2490389e+33 * -1.4242695e-17 = 3.2032375e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000100000001100000101101110100;
		b = 32'b10111110011010100000101011011101;
		correct = 32'b00000010111101010001100001010000;
		#400 //-1.5756883e-36 * -0.22855707 = 3.601347e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100010010010011001100001000001;
		b = 32'b10110010110011111000101001000110;
		correct = 32'b11010101101000110110111100000000;
		#400 //9.2969165e+20 * -2.4160851e-08 = -22462142000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011111111111110111010011110111;
		b = 32'b01001110111001110111000000011101;
		correct = 32'b10101111011001101111001001101011;
		#400 //-1.081902e-19 * 1941442200.0 = -2.1004502e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100001101111100011110100011011;
		b = 32'b10010001101111011011011101010111;
		correct = 32'b10110100000011001111101101011011;
		#400 //4.3866056e+20 * -2.9931934e-28 = -1.3129959e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111110110001000111101000110101;
		b = 32'b01000110000111110110100101011011;
		correct = 32'b11000101011101001011000110000110;
		#400 //-0.38374487 * 10202.339 = -3915.0952
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110011110100111101110001110101;
		b = 32'b11110100111000011010010000111000;
		correct = 32'b11101001001110101011110010101010;
		#400 //9.865554e-08 * -1.4301728e+32 = -1.4109446e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010011000000110101110101100;
		b = 32'b01001111100100101011001100010011;
		correct = 32'b11001010100000001001101001100100;
		#400 //-0.0008560966 * 4922418700.0 = -4214066.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011101110110111011011110011011;
		b = 32'b11000000001100110010000111011111;
		correct = 32'b00011110100110011011111001110011;
		#400 //-5.815866e-21 * -2.7989423 = 1.6278273e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100001101101001000000011000000;
		b = 32'b11011100101111110001111111010110;
		correct = 32'b01111111000001101100001010000010;
		#400 //-4.1621142e+20 * -4.303738e+17 = 1.791265e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010000100100010001111000010001;
		b = 32'b11010011100010100000111010010010;
		correct = 32'b00100100100111001000010011101111;
		#400 //-5.723874e-29 * -1185899900000.0 = 6.7879414e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100010001101100101001111100110;
		b = 32'b10011010111000011110110011000101;
		correct = 32'b10111101101000001110100001011111;
		#400 //8.4083824e+20 * -9.344034e-23 = -0.07856821
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110111011011000111111001101110;
		b = 32'b10000000100100101101100000111101;
		correct = 32'b10111000100001111010011111011110;
		#400 //4.7966655e+33 * -1.3485554e-38 = -6.468569e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100010010011111011010111100101;
		b = 32'b01110000001010101011110011001100;
		correct = 32'b11010011000010101000011111111001;
		#400 //-2.8150025e-18 * 2.1136277e+29 = -594986700000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010111000000101000001100001010;
		b = 32'b00100011100101011000100001001011;
		correct = 32'b10111011000110000111011110000001;
		#400 //-143499320000000.0 * 1.6212335e-17 = -0.002326459
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011111000111100010111111111100;
		b = 32'b01000011001001001011101100000011;
		correct = 32'b01100010110010111001010010011001;
		#400 //1.1398606e+19 * 164.73051 = 1.8776983e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111111110010010000110011101100;
		b = 32'b00010011010100010011110110110011;
		correct = 32'b10010011101001000101010000000001;
		#400 //-1.5707068 * 2.6409929e-27 = -4.1482255e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111011100001101110100101011111;
		b = 32'b00010100010010001001001001000110;
		correct = 32'b00010000010100110110011011010000;
		#400 //0.0041171755 * 1.0126267e-26 = 4.1691617e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000000101001000101100000011;
		b = 32'b11000001010100101010101011001101;
		correct = 32'b00110001111101000111101001000111;
		#400 //-5.4039634e-10 * -13.166699 = 7.115236e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111101000100010101011111101011;
		b = 32'b10111101001110010011001110111101;
		correct = 32'b10111010110100100100101111010001;
		#400 //0.035484236 * -0.045215357 = -0.0016044324
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010101110010010101110100101001;
		b = 32'b00101100101101011101010010001101;
		correct = 32'b00000011000011110000011000001110;
		#400 //8.1330234e-26 * 5.1679273e-12 = 4.2030873e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110001101010101010001101101110;
		b = 32'b10011101101100100100110101111001;
		correct = 32'b11001111111011011011001010001101;
		#400 //1.6899208e+30 * -4.7196313e-21 = -7975803400.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001110101111101100000101100001;
		b = 32'b00101111100001001011001111011001;
		correct = 32'b00111110110001011100001101110010;
		#400 //1600172200.0 * 2.413845e-10 = 0.38625675
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011011111101110010010100000010;
		b = 32'b11100110100010100011000110010000;
		correct = 32'b11000011000001010110100111001100;
		#400 //4.0886638e-22 * -3.2630042e+23 = -133.41327
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111001111100101110101101010101;
		b = 32'b11101101101000011111111111100000;
		correct = 32'b01101000000110011011100011001101;
		#400 //-0.00046333173 * -6.2670526e+27 = 2.9037242e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000010110000100110100110011010;
		b = 32'b11010010101001110101111100011011;
		correct = 32'b00010101111111100011011000111010;
		#400 //-2.856635e-37 * -359427570000.0 = 1.0267534e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101011001000111110111101101000;
		b = 32'b00011101111111111111010100110111;
		correct = 32'b10001001101000111110100010000000;
		#400 //-5.8241476e-13 * 6.7751484e-21 = -3.9459465e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111000111010111011010010110100;
		b = 32'b01111000001000011010000011101011;
		correct = 32'b11110001100101001101000011001111;
		#400 //-0.00011239332 * 1.3112869e+34 = -1.4737989e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000000101100110100011110101101;
		b = 32'b11101011010010010101000010111000;
		correct = 32'b00101100100011001111101111001110;
		#400 //-1.6464266e-38 * -2.4337527e+26 = 4.0069953e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001111101101100101100110110111;
		b = 32'b01110111010010000111111110000111;
		correct = 32'b11000111100011101101000011101110;
		#400 //-1.7981142e-29 * 4.0665857e+33 = -73121.86
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110011111110000111101110001101;
		b = 32'b10001100110011010010000111011011;
		correct = 32'b01000001010001110001101111001100;
		#400 //-3.9373643e+31 * -3.1605627e-31 = 12.444286
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101011000111011101000111111010;
		b = 32'b10110100101100111111011111011110;
		correct = 32'b00100000010111011110010101000001;
		#400 //-5.6069006e-13 * -3.3521695e-07 = 1.8795282e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000010001100110100111011110111;
		b = 32'b11100111111011011001110111011111;
		correct = 32'b01101010101001100110111010101110;
		#400 //-44.827114 * -2.2442261e+24 = 1.0060218e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111011010001100000101000111100;
		b = 32'b10010110110000110001011110001010;
		correct = 32'b01010010100101101110110000000001;
		#400 //-1.02828236e+36 * -3.1518804e-25 = 324102300000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100011001001111001101100000001;
		b = 32'b11110100110101011101101111111101;
		correct = 32'b01011000100011000000001111111111;
		#400 //-9.0859115e-18 * -1.3554945e+32 = 1231590300000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111100001010001110100001111101;
		b = 32'b01100110010110011101000100111001;
		correct = 32'b01100011000011111011011100011101;
		#400 //0.010309336 * 2.5715325e+23 = 2.651079e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001011101000111000100001001011;
		b = 32'b11010101100101001010011100000111;
		correct = 32'b00100001101111011110101011111011;
		#400 //-6.2990387e-32 * -20430637000000.0 = 1.2869337e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001111010111000111010001001011;
		b = 32'b00010000001010110111111010000110;
		correct = 32'b00100000000100111010111010100011;
		#400 //3698609000.0 * 3.3821274e-29 = 1.2509167e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100100101010110010101000101000;
		b = 32'b00010111010000011000001100111100;
		correct = 32'b00111100100000010110001010000111;
		#400 //2.5259447e+22 * 6.2527304e-25 = 0.015794052
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101100111001000110111001010000;
		b = 32'b00011001100110101100110001100000;
		correct = 32'b11000111000010100010000010111010;
		#400 //-2.2092482e+27 * 1.6005773e-23 = -35360.727
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100111000100110010000000000110;
		b = 32'b00100111111110010111101001010010;
		correct = 32'b10001111100011110110000001110010;
		#400 //-2.0417708e-15 * 6.9244003e-15 = -1.4138038e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101110001111111010011100111010;
		b = 32'b00111000000100001000110100111000;
		correct = 32'b01100110110110000110111110010011;
		#400 //1.482845e+28 * 3.4463796e-05 = 5.1104467e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011101111101110101101111111010;
		b = 32'b00000010100101010010011111111010;
		correct = 32'b10100001000100000001111100101001;
		#400 //-2.2280144e+18 * 2.1916528e-37 = -4.883034e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010001111001010101100101101000;
		b = 32'b01101011100111001010011110111000;
		correct = 32'b00111110000011000101100010111110;
		#400 //3.618493e-28 * 3.787689e+26 = 0.13705727
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000001100001101000011111100101;
		b = 32'b01000011000110001101001100100110;
		correct = 32'b00000101001000001001111101001100;
		#400 //4.9418825e-38 * 152.8248 = 7.552422e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011111101101110001011000000001;
		b = 32'b01011110010111100101000010010110;
		correct = 32'b10111110100111101111111010110111;
		#400 //-7.753992e-20 * 4.0048672e+18 = -0.31053707
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010100000100111101100001101;
		b = 32'b00111001010001001000011100100111;
		correct = 32'b10110100010010000101011000110001;
		#400 //-0.0009954885 * 0.00018742365 = -1.8657808e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010000001000100111100011000010;
		b = 32'b10000110101110111111000100111010;
		correct = 32'b00010111011011101000111010011100;
		#400 //-10903292000.0 * -7.069603e-35 = 7.7081946e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111101000011011100001110111010;
		b = 32'b01100001100000111101000000010101;
		correct = 32'b11011111000100011111110011000110;
		#400 //-0.034610488 * 3.0393967e+20 = -1.05195e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010011000100011000001011111110;
		b = 32'b11011001101001101001101110100110;
		correct = 32'b01101101001111010110011011010011;
		#400 //-624967940000.0 * -5861998000000000.0 = 3.663561e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100101101110100011110010000000;
		b = 32'b00110111101000110011010110000010;
		correct = 32'b10011101111011010111011011100101;
		#400 //-3.2306853e-16 * 1.945603e-05 = -6.285631e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001011010101001111011100001100;
		b = 32'b10111101101000101001011100011101;
		correct = 32'b00001001100001110100001000001011;
		#400 //-4.1015572e-32 * -0.07938979 = 3.2562174e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110111000111111010011100101;
		b = 32'b11100111010001110111010101111101;
		correct = 32'b01011110101100011001101111111100;
		#400 //-6.7936367e-06 * -9.419182e+23 = 6.39905e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000010001110010100011101101010;
		b = 32'b10101100100000110111110011011100;
		correct = 32'b10101111001111100101001111010010;
		#400 //46.31974 * -3.737106e-12 = -1.7310178e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101111010010000001111110111001;
		b = 32'b01101010001100100001010110000001;
		correct = 32'b11011010000010110011011011011110;
		#400 //-1.8201164e-10 * 5.3822586e+25 = -9796337000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101110110110010111011010011110;
		b = 32'b00010000011110011000011011010101;
		correct = 32'b00111111110100111111011011101001;
		#400 //3.3650823e+28 * 4.9210462e-29 = 1.6559726
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110010010011100101011011111010;
		b = 32'b11110010101000101100100110000010;
		correct = 32'b01100101100000110011010101110101;
		#400 //-1.2010554e-08 * -6.448663e+30 = 7.7452015e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101101001100011110100110111101;
		b = 32'b11000100110111001011001010010001;
		correct = 32'b01110010100110010110000011111000;
		#400 //-3.4413387e+27 * -1765.5802 = 6.0759596e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011010001001101011101101100001;
		b = 32'b01001010100010010000101101101011;
		correct = 32'b11100101001100101000001101101101;
		#400 //-1.1732718e+16 * 4490677.5 = -5.268785e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010110101101010110011001110101;
		b = 32'b11110011001100111010011111101101;
		correct = 32'b01001010011111101001101101000011;
		#400 //-2.9306787e-25 * -1.4233812e+31 = 4171472.8
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001110101000111111011010010111;
		b = 32'b00111011001111011011101110010001;
		correct = 32'b01001010011100110000101001011111;
		#400 //1375423400.0 * 0.002895091 = 3981975.8
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100111010010001110111001101111;
		b = 32'b00110000111100010010000101001001;
		correct = 32'b00011000101111010100001010010111;
		#400 //2.788483e-15 * 1.7544518e-09 = 4.8922593e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110010000011100100101001001010;
		b = 32'b00001011000010110011111001100101;
		correct = 32'b00111101100110101100101000001001;
		#400 //2.8183476e+30 * 2.6817367e-32 = 0.075580664
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101101110101110101010000101100;
		b = 32'b01001101010010011011001010001111;
		correct = 32'b10111011101010011010011101000111;
		#400 //-2.448005e-11 * 211495150.0 = -0.0051774117
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111001001001011001011011100000;
		b = 32'b11011111001111000011110001100001;
		correct = 32'b01011000111100111000001110110101;
		#400 //-0.00015791832 * -1.3563823e+19 = 2141976000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101100001001110110111010110100;
		b = 32'b10011110011000101101000010011010;
		correct = 32'b00001011000101000101100000101010;
		#400 //-2.379358e-12 * -1.2007478e-20 = 2.857009e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000011001001110100011111101000;
		b = 32'b01001011111000011110011001101100;
		correct = 32'b10001111100100111001110011000100;
		#400 //-4.9159433e-37 * 29609176.0 = -1.4555703e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011010110100101010110011111110;
		b = 32'b00110100101101100100110001000001;
		correct = 32'b01010000000101100000010110111101;
		#400 //2.9649976e+16 * 3.3955624e-07 = 10067834000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101111000111010010010101101001;
		b = 32'b00011111101001000010110001010101;
		correct = 32'b00001111010010011000111001011100;
		#400 //1.4292358e-10 * 6.953004e-20 = 9.9374825e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110000100000100101111101010;
		b = 32'b10111100000011011101100100110011;
		correct = 32'b00110010100111111110100001111010;
		#400 //-2.150186e-06 * -0.008657741 = 1.8615754e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101010101100010111110010101101;
		b = 32'b10101011010001001010000011111001;
		correct = 32'b00010110100010000101001100001111;
		#400 //-3.1528027e-13 * -6.985658e-13 = 2.2024402e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111100000000100010010101000011;
		b = 32'b11110010000101000111001010111010;
		correct = 32'b01101110100101101110111110111100;
		#400 //-0.007943454 * -2.9403186e+30 = 2.3356286e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011011000101110111001100100010;
		b = 32'b11011101011110100000100101111010;
		correct = 32'b10111001000100111110110000001010;
		#400 //1.2527629e-22 * -1.1260666e+18 = -0.00014106944
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100100100000111010100111110001;
		b = 32'b01001000110100000010100011001010;
		correct = 32'b00101101110101100001111000011101;
		#400 //5.7100086e-17 * 426310.3 = 2.4342356e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010100111101110111100101111000;
		b = 32'b10110000100001111010010111110011;
		correct = 32'b01000110000000110010000101111010;
		#400 //-8503158600000.0 * -9.869708e-10 = 8392.369
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011010001010111100011000110011;
		b = 32'b10111100110101111010101011010011;
		correct = 32'b10010111100100001011011000010100;
		#400 //3.5522075e-23 * -0.026326573 = -9.351745e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101101111000000111001110011100;
		b = 32'b11110010000101101011010010000110;
		correct = 32'b11100000100001000010001000000100;
		#400 //2.5517193e-11 * -2.9850234e+30 = -7.616942e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001111010110011100001000101101;
		b = 32'b11010111100000111110101010010110;
		correct = 32'b11100111011000000110101111010000;
		#400 //3653381400.0 * -290087120000000.0 = -1.0597989e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010101100100001110010000011011;
		b = 32'b00111101110111000100110001000000;
		correct = 32'b01010011111110010101111001011110;
		#400 //19913672000000.0 * 0.10756731 = 2142060200000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001100100101100000001101011001;
		b = 32'b00111000101000111100110101011110;
		correct = 32'b10000101101111111111100011110011;
		#400 //-2.3113174e-31 * 7.810698e-05 = -1.8053003e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011000010101010100100110100101;
		b = 32'b00101000111001000001101111110100;
		correct = 32'b10000001101111100000110011100001;
		#400 //-2.7566786e-24 * 2.5325208e-14 = -6.981346e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110100101110000111101100000100;
		b = 32'b01110011000011101101001110111111;
		correct = 32'b11101000010011011101100110100111;
		#400 //-3.4362176e-07 * 1.1315931e+31 = -3.8884004e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010010001001110111010001100111;
		b = 32'b10100110010100111100010000110111;
		correct = 32'b00111001000010101000010101001010;
		#400 //-179803110000.0 * -7.347125e-16 = 0.0001321036
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010101011110111101110011100101;
		b = 32'b11100100010011011100110011001111;
		correct = 32'b11111010010010100111100101100011;
		#400 //17307885000000.0 * -1.5185362e+22 = -2.628265e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011011001111111000000000010101;
		b = 32'b01100001101010111101111111100001;
		correct = 32'b00111101100000001001001000000111;
		#400 //1.5840535e-22 * 3.9631568e+20 = 0.062778525
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100101101011000001000001100100;
		b = 32'b10110100000110111001010111001010;
		correct = 32'b01011010010100010010010100110100;
		#400 //-1.0156867e+23 * -1.4489993e-07 = 1.4717294e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000010110011110111110011110110;
		b = 32'b00001010101000111101101100011110;
		correct = 32'b00001110000001001100111000101001;
		#400 //103.744064 * 1.5778752e-32 = 1.6369519e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100100000001101111000000011100;
		b = 32'b01100101100111110000101100101101;
		correct = 32'b11001010001001111010101000001011;
		#400 //-2.926e-17 * 9.38828e+22 = -2747010.8
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100000000101100001011010010010;
		b = 32'b10100000011111111110011000101000;
		correct = 32'b01000001000101100000011101101011;
		#400 //-4.325997e+19 * -2.1675492e-19 = 9.376811
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110001111100100100000010000000;
		b = 32'b10111000100101000011001110000110;
		correct = 32'b10101011000011000011111000001100;
		#400 //7.0504598e-09 * -7.066787e-05 = -4.98241e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100111000101111100011001101101;
		b = 32'b10000101100000110010011100100000;
		correct = 32'b00101101000110111000001101111000;
		#400 //-7.1673765e+23 * -1.2333553e-35 = 8.839922e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100101010111000011101011111;
		b = 32'b01000101011101011111011011110101;
		correct = 32'b01001010101001001100111000000110;
		#400 //1372.2303 * 3935.4348 = 5400323.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101110111101110001010010000110;
		b = 32'b11101111110010101011111001101101;
		correct = 32'b01011111010000111010110111111100;
		#400 //-1.1235905e-10 * -1.25492365e+29 = 1.4100203e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010110000100110010001111101001;
		b = 32'b01010011000101101000100101010010;
		correct = 32'b11101001101011010000101111110000;
		#400 //-40445610000000.0 * 646548950000.0 = -2.6150068e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100110101000000011010000101100;
		b = 32'b00100001110001010010100000101100;
		correct = 32'b01001000111101101100001010010011;
		#400 //3.7827052e+23 * 1.3359873e-18 = 505364.6
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100111100101100111111100001111;
		b = 32'b11010111000100100011101111111000;
		correct = 32'b01111111001010111110111101101111;
		#400 //-1.4213976e+24 * -160786260000000.0 = 2.285412e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000100101101100100010101000101;
		b = 32'b00000000001100010000110011000010;
		correct = 32'b10000101000010111011000101011110;
		#400 //-1458.1647 * 4.504516e-39 = -6.568326e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110100101000110111001100011100;
		b = 32'b11100110011001110100011000100111;
		correct = 32'b01011011100100111010100110101001;
		#400 //-3.044487e-07 * -2.7304018e+23 = 8.312673e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111111001110010000110100101000;
		b = 32'b00011111110100100000101001111000;
		correct = 32'b10011111100101111101010001011100;
		#400 //-0.722857 * 8.895578e-20 = -6.4302307e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000011110111010100011100011001;
		b = 32'b11110100010101011010110010001011;
		correct = 32'b01111000101110001011000101001100;
		#400 //-442.55545 * -6.771599e+31 = 2.9968082e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010110101110000010000100000011;
		b = 32'b10000010100010100000010100001011;
		correct = 32'b00011001110001101000101011011000;
		#400 //-101225960000000.0 * -2.0280172e-37 = 2.0528799e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111001110011110100101001011000;
		b = 32'b11101101101110110001011010000100;
		correct = 32'b01101000000101110111110110001010;
		#400 //-0.00039537507 * -7.2376146e+27 = 2.8615725e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100000000001111100111100101100;
		b = 32'b10100001110110000001000001011001;
		correct = 32'b01000010011001010011111011110011;
		#400 //-3.9144356e+19 * -1.4641057e-18 = 57.311474
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101101011010000101110001010101;
		b = 32'b00101001011110010110001111001010;
		correct = 32'b11010111011000100101110001100010;
		#400 //-4.494509e+27 * 5.537566e-14 = -248886410000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101011100111000011000000011010;
		b = 32'b10001011010011000011010011000110;
		correct = 32'b00110111011110010010110100001111;
		#400 //-3.7763916e+26 * -3.9328673e-32 = 1.4852048e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100100001101010011100111010011;
		b = 32'b01101100110110100111110010011000;
		correct = 32'b11010001100110101010101101110001;
		#400 //-3.9297098e-17 * 2.1130736e+27 = -83037660000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110111100100111000110101000111;
		b = 32'b11111001110100101110110100100111;
		correct = 32'b11110001111100110010010100101001;
		#400 //1.7589553e-05 * -1.3689905e+35 = -2.407993e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001010100010000000000101111000;
		b = 32'b11010001011110001101000100000110;
		correct = 32'b00011100100001000011000001111001;
		#400 //-1.3096876e-32 * -66791170000.0 = 8.747557e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111100110010001010011011100010;
		b = 32'b00001110101111100000010000010010;
		correct = 32'b11001100000101001110111100001100;
		#400 //-8.334753e+36 * 4.6842536e-30 = -39042096.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100111100100001000000111110010;
		b = 32'b00101100010101111001011100011001;
		correct = 32'b01010100011100110110010011011010;
		#400 //1.3648357e+24 * 3.0637214e-12 = 4181476200000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000011111011001010000100101000;
		b = 32'b10000111101100001001010100100010;
		correct = 32'b00001100001000110011100010100101;
		#400 //-473.25903 * -2.656919e-34 = 1.2574109e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000101110010100100010010110010;
		b = 32'b01100100100011111110010001000101;
		correct = 32'b01101010111000110110000101110110;
		#400 //6472.587 * 2.1234664e+22 = 1.374432e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001010010001111101101000101100;
		b = 32'b10011000011110101110010000110111;
		correct = 32'b00100011010000111101110100111000;
		#400 //-3274379.0 * -3.2426962e-24 = 1.0617816e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101111111110010011100101111100;
		b = 32'b10010101010111011001110011001011;
		correct = 32'b00000101110101111011111101000101;
		#400 //-4.533368e-10 * -4.4754282e-26 = 2.0288764e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101111111001010110001000100001;
		b = 32'b01101111110000000001011011111100;
		correct = 32'b11100000001011000001111000110001;
		#400 //-4.1724582e-10 * 1.1889782e+29 = -4.9609617e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100011010001000100010101101010;
		b = 32'b11010111110001110101010010011000;
		correct = 32'b10111011100110001101001011010001;
		#400 //1.063988e-17 * -438332280000000.0 = -0.004663803
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001101011000000101000111010001;
		b = 32'b00111001011000011010110111111101;
		correct = 32'b11000111010001011100000001011110;
		#400 //-235216140.0 * 0.00021522488 = -50624.367
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111011110011101110110110100000;
		b = 32'b10011101001010010001111110101111;
		correct = 32'b11011001100010001011010001111011;
		#400 //2.1488655e+36 * -2.2383344e-21 = -4809879700000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110101010011111100010001101101;
		b = 32'b00001111101100111000000110110011;
		correct = 32'b11000101100100011010111110011011;
		#400 //-2.6337633e+32 * 1.7700721e-29 = -4661.9507
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110100001100110100010001110111;
		b = 32'b10010111101000001010110010110110;
		correct = 32'b01001100011000010000011101111000;
		#400 //-5.681212e+31 * -1.0383356e-24 = 58990050.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110101101010001110000000110111;
		b = 32'b11001111101101110101101011110111;
		correct = 32'b11000101111100011110100010010010;
		#400 //1.258223e-06 * -6152384000.0 = -7741.0713
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111001001010000010111000110010;
		b = 32'b00011100001000001100111101000000;
		correct = 32'b11010101110100110100101000001101;
		#400 //-5.4577677e+34 * 5.3207424e-22 = -29039375000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000011010001001001000011001111;
		b = 32'b01010110111001101000101110100101;
		correct = 32'b00011010101100010000010101010011;
		#400 //5.7765455e-37 * 126743720000000.0 = 7.3214086e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001101011101010100010001100010;
		b = 32'b10111110010101000111000011100000;
		correct = 32'b11001100010010111000100011000110;
		#400 //257181220.0 * -0.20746183 = -53355290.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110000110100111011010111100001;
		b = 32'b10010101010101110000110100101110;
		correct = 32'b10000110101100011101100010100110;
		#400 //1.5403964e-09 * -4.34293e-26 = -6.6898336e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101101010100010101110101101101;
		b = 32'b10001010111100011011111100110011;
		correct = 32'b10111000110001011011010101010010;
		#400 //4.049707e+27 * -2.3279377e-32 = -9.4274656e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001001000110110001111001111111;
		b = 32'b01001011101101000110100101100110;
		correct = 32'b10010101010110101010001010011101;
		#400 //-1.8671786e-33 * 23646924.0 = -4.415303e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010001010110000000011100110000;
		b = 32'b00110001010100001000101111101011;
		correct = 32'b01000011001011111111101111101001;
		#400 //57989595000.0 * 3.0347518e-09 = 175.98402
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100000001011111000110111111001;
		b = 32'b00111001111100001101100000111110;
		correct = 32'b10011010101001010010100101100100;
		#400 //-1.4870051e-19 * 0.0004593748 = -6.830927e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010111000101011011110110001101;
		b = 32'b01000011110010010101101000101101;
		correct = 32'b00011011011010111000110100100101;
		#400 //4.8383743e-25 * 402.7045 = 1.9484351e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111011001010110001000011110010;
		b = 32'b00011100111001101110110011000100;
		correct = 32'b00011000100110100100111101110000;
		#400 //0.002610263 * 1.5281326e-21 = 3.988828e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000101110111000101011101111110;
		b = 32'b01101110100111111000001110110101;
		correct = 32'b11110101000010010100101110110100;
		#400 //-7050.9365 * 2.468367e+28 = -1.74043e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001100011100111110000000110110;
		b = 32'b00000000001010111010110001100110;
		correct = 32'b10001100101001100110101110010100;
		#400 //-63930584.0 * 4.010771e-39 = -2.5641096e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010011010010100001100000011101;
		b = 32'b01001100010101000011100000101111;
		correct = 32'b10100000001001111000100001010010;
		#400 //-2.5507873e-27 * 55632060.0 = -1.4190555e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111001111001101001011011011111;
		b = 32'b11001001111010000100101110011001;
		correct = 32'b01000100010100010011110011010010;
		#400 //-0.00043981426 * -1902963.1 = 836.9503
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011011100001001001111111011100;
		b = 32'b01101000010101111011100110001011;
		correct = 32'b11000100010111111000010011000011;
		#400 //-2.1940875e-22 * 4.0749258e+24 = -894.0744
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001100000010001011111000100011;
		b = 32'b00000010111100000100011100111001;
		correct = 32'b00001111100000000101100001001100;
		#400 //35846284.0 * 3.530571e-37 = 1.2655785e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100010100000100011111111111010;
		b = 32'b11001010011101101011000110000010;
		correct = 32'b01101101011110110000011110010101;
		#400 //-1.2013434e+21 * -4041824.5 = 4.855619e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110010001110110111011111101100;
		b = 32'b01000000111100000011010011010111;
		correct = 32'b11110011101011111110011100011111;
		#400 //-3.713195e+30 * 7.50645 = -2.7872914e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010001111110000110011101110000;
		b = 32'b00101000110011010011101110011010;
		correct = 32'b00111011010001110010010010101010;
		#400 //133360910000.0 * 2.278542e-14 = 0.0030386844
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100101000110010111000110011000;
		b = 32'b00101001001100000101101100100000;
		correct = 32'b01001110110100110110100101101110;
		#400 //4.5288594e+22 * 3.915889e-14 = 1773451000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011100000101110001001001000100;
		b = 32'b10100000110110011101011100101010;
		correct = 32'b10111101100000001000110101110101;
		#400 //1.7009122e+17 * -3.6903614e-19 = -0.06276981
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111101111011110011010000101101;
		b = 32'b00001100011011010000000001010001;
		correct = 32'b00001010110111010111001110011001;
		#400 //0.116798736 * 1.8257911e-31 = 2.1325009e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011111110011110110001011100110;
		b = 32'b10101100110011110101010000000100;
		correct = 32'b00001101001001111111010100001000;
		#400 //-8.7831524e-20 * -5.8926215e-12 = 5.1755794e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110011000111000000110000001101;
		b = 32'b10101101101100000110010100100110;
		correct = 32'b10100001010101110000101111100010;
		#400 //3.633254e-08 * -2.0053802e-11 = -7.286056e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110010111011101100111111101000;
		b = 32'b11001011011011100000100011110001;
		correct = 32'b10111110110111100000110110100001;
		#400 //2.7801391e-08 * -15599857.0 = -0.43369773
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100011110011001001111101101100;
		b = 32'b01001000001010000011011001111101;
		correct = 32'b10101100100001100111010000101100;
		#400 //-2.2185242e-17 * 172249.95 = -3.8214067e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000011011100110000101110001001;
		b = 32'b11101100000000101111110111100010;
		correct = 32'b00101111111110001011100111001001;
		#400 //-7.1424524e-37 * -6.3343714e+26 = 4.5242946e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011011100100001100011001000101;
		b = 32'b10101100110001110010001101110101;
		correct = 32'b10001000111000010011110001011010;
		#400 //2.395093e-22 * -5.6598567e-12 = -1.35558835e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101010001000011010110110101010;
		b = 32'b10110011100101001000111100100111;
		correct = 32'b10011110001110111010010110011110;
		#400 //1.4359924e-13 * -6.917826e-08 = -9.933946e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110101101110101100100100011100;
		b = 32'b10010011011001010010111111000101;
		correct = 32'b10001001101001110011100011000001;
		#400 //1.391661e-06 * -2.8927416e-27 = -4.025716e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000101111001000011000010111101;
		b = 32'b00100001100010101000100111001010;
		correct = 32'b00100111111101101111101000110000;
		#400 //7302.0923 * 9.387716e-19 = 6.854997e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111100010010111111111001110111;
		b = 32'b01100110101001011010000111101000;
		correct = 32'b01100011100000111111110000000111;
		#400 //0.012450806 * 3.9108856e+23 = 4.869368e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011010010001110101110100010;
		b = 32'b01011110010101111000100110011011;
		correct = 32'b11101010001010010010100111100101;
		#400 //-13167522.0 * 3.8827788e+18 = -5.1126576e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000101110110100010101100010101;
		b = 32'b11111011001011101011000101111011;
		correct = 32'b01000001100101001110000010001001;
		#400 //-2.0516447e-35 * -9.070594e+35 = 18.609636
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110010110110000001100010010010;
		b = 32'b11000110010110110111111011000101;
		correct = 32'b10111001101110010100100000000111;
		#400 //2.5156883e-08 * -14047.692 = -0.00035339614
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011001100000110001000100110010;
		b = 32'b11100111011100110001110000110110;
		correct = 32'b01000001011110001110111110001000;
		#400 //-1.3552028e-23 * -1.14805546e+24 = 15.558479
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011000001100000100111010111001;
		b = 32'b01101101001111110101010010101000;
		correct = 32'b01000110000000111100010100001010;
		#400 //2.2787212e-24 * 3.7008738e+27 = 8433.26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101010010100101001001100110011;
		b = 32'b10101000110011110001011101100000;
		correct = 32'b01010011101010100101100001000000;
		#400 //-6.3642388e+25 * -2.2991754e-14 = 1463250000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010100000010101011101101101011;
		b = 32'b10010101110110100001001101100011;
		correct = 32'b10101010011011000101110000110101;
		#400 //2383399400000.0 * -8.8080086e-26 = -2.0993001e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101000011010111000010010011101;
		b = 32'b00101100010100101011101101110011;
		correct = 32'b01010101010000011101111100111100;
		#400 //4.4488096e+24 * 2.994685e-12 = 13322783000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111000000001110101010101000100;
		b = 32'b10100011001111100110111000010110;
		correct = 32'b10011011110010010101011011110101;
		#400 //3.2265918e-05 * -1.0323232e-17 = -3.3308855e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100000101110110111110101001010;
		b = 32'b01111101001010100000101001001010;
		correct = 32'b11011110011110010001000101111000;
		#400 //-3.1761942e-19 * 1.4126386e+37 = -4.4868145e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011010011100100110010000111011;
		b = 32'b11010100110010000000110100101111;
		correct = 32'b00101111101111010110101011001010;
		#400 //-5.0125393e-23 * -6873717000000.0 = 3.4454778e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111011001110010100100110001000;
		b = 32'b10101011000010000001110110101111;
		correct = 32'b10100110110001010000100100011000;
		#400 //0.0028272588 * -4.83581e-13 = -1.3672086e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110100101101101111101000000111;
		b = 32'b10100011011101101011010010100001;
		correct = 32'b00011000101100000101010101011110;
		#400 //-3.408206e-07 * -1.3373936e-17 = 4.5581133e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111000010111001111101111010111;
		b = 32'b11111110000101110110011111100100;
		correct = 32'b01110111000000101011001000111010;
		#400 //-5.268663e-05 * -5.0313215e+37 = 2.6508338e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011111101010110011110000000110;
		b = 32'b00010111000100011100010111110110;
		correct = 32'b00110111010000110000001011010010;
		#400 //2.4677487e+19 * 4.710189e-25 = 1.1623562e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101010110100001001011100010110;
		b = 32'b11011010101100100110010110011110;
		correct = 32'b01000110000100010101101111011010;
		#400 //-3.705306e-13 * -2.5107138e+16 = 9302.963
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111100000000110001001010000111;
		b = 32'b10010011011101000111011111011100;
		correct = 32'b10001111111110100101011000001110;
		#400 //0.008000023 * -3.0856225e-27 = -2.468505e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000000000100111001001101100110;
		b = 32'b01111110010101000000000100000001;
		correct = 32'b00111110000000011011000100100001;
		#400 //1.797751e-39 * 7.0450387e+37 = 0.12665226
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010100001101000101100000101011;
		b = 32'b10110111111101011110100101101101;
		correct = 32'b01001100101011010011110011010010;
		#400 //-3098293300000.0 * -2.9314973e-05 = 90826380.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010110001100010111110110100110;
		b = 32'b00000000001101000101000110010000;
		correct = 32'b00010110100100010001100001001001;
		#400 //48788304000000.0 * 4.804705e-39 = 2.344134e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001111111100010100000110001111;
		b = 32'b11100110110100010000110000001101;
		correct = 32'b11110111010001010000000111100001;
		#400 //8095211000.0 * -4.9359845e+23 = -3.9957836e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010010111110101101001100100011;
		b = 32'b11000001101100000111100001000101;
		correct = 32'b10010101001011001110011011111111;
		#400 //1.5829267e-27 * -22.058725 = -3.4917347e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011110100100110100110011000111;
		b = 32'b11000101111010000101001010101101;
		correct = 32'b00100101000001011010110100100110;
		#400 //-1.5595985e-20 * -7434.3345 = 1.1594576e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010001011001001101111111001011;
		b = 32'b11100101101000111110101101010111;
		correct = 32'b10110111100100101000110011100101;
		#400 //1.805499e-28 * -9.676087e+22 = -1.7470165e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001101001110010010110111001111;
		b = 32'b00110011001110001011110010011010;
		correct = 32'b10000001000001011010000101011010;
		#400 //-5.7062666e-31 * 4.301237e-08 = -2.4544006e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101011000100101100101111000001;
		b = 32'b00111011001001000000101001001110;
		correct = 32'b01100110101111000010000011100001;
		#400 //1.7746537e+26 * 0.0025030556 = 4.442057e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110010010011101011000101011010;
		b = 32'b10111101111100110111111110010001;
		correct = 32'b01110000110001001001100101010111;
		#400 //-4.0939723e+30 * -0.11889566 = 4.867555e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001110011100011000010010000001;
		b = 32'b01100101001000000101010001010000;
		correct = 32'b01110100000101110100001001011100;
		#400 //1012998200.0 * 4.732087e+22 = 4.793596e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101101100010100111000110000010;
		b = 32'b11010010011111000111111111100000;
		correct = 32'b11000000100010001000110011100011;
		#400 //1.5739191e-11 * -271119290000.0 = -4.267198
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100100000110111100011000111010;
		b = 32'b10100110011101011100100100101100;
		correct = 32'b01001011000101011000111100011111;
		#400 //-1.1494116e+22 * -8.527409e-16 = 9801503.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100000011000001000111001011001;
		b = 32'b01001100001111010101010011101111;
		correct = 32'b00101101001001100001001110011000;
		#400 //1.9020637e-19 * 49632188.0 = 9.440358e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011011101001001011100011000110;
		b = 32'b00101110000110010001111011000111;
		correct = 32'b00001010010001010000110001111000;
		#400 //2.725093e-22 * 3.4815508e-11 = 9.48755e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110010100101001010110000100110;
		b = 32'b11101010101001101101100101011001;
		correct = 32'b11011101110000011100101110110101;
		#400 //1.7307752e-08 * -1.0085404e+26 = -1.7455568e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110000101110001100110111000111;
		b = 32'b01011001100110111001011100010001;
		correct = 32'b01001010111000001010001101001010;
		#400 //1.3446247e-09 * 5474340000000000.0 = 7360933.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000011101110001001101110110100;
		b = 32'b00101000011101011101110100100001;
		correct = 32'b10101100101100010100110001111001;
		#400 //-369.21643 * 1.3648182e-14 = -5.0391327e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000110101101111100001001110100;
		b = 32'b10100011101000000100001000111110;
		correct = 32'b10101010111001100001001000101010;
		#400 //23521.227 * -1.737529e-17 = -4.086881e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100111110100000101110100000101;
		b = 32'b10100111101101011001100010110111;
		correct = 32'b00010000000100111100111000010001;
		#400 //-5.783245e-15 * -5.0403166e-15 = 2.9149386e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010110010100110011100110101101;
		b = 32'b00010011010110110111100011000100;
		correct = 32'b00101010001101010001010111111100;
		#400 //58061167000000.0 * 2.7701228e-27 = 1.6083657e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101100111101110111111100000000;
		b = 32'b10010111110000010101110001111111;
		correct = 32'b01000101001110101111000000101011;
		#400 //-2.3936353e+27 * -1.2495682e-24 = 2991.0105
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110001010110010011010110111110;
		b = 32'b01111101101001111101001011111100;
		correct = 32'b11101111100011100110010100010011;
		#400 //-3.1608205e-09 * 2.788457e+37 = -8.8138125e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011111101101000011001001001001;
		b = 32'b01000111111111101101011000000000;
		correct = 32'b00101000001100110110000010000110;
		#400 //7.6316155e-20 * 130476.0 = 9.957426e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011000010111101101101011101010;
		b = 32'b10011001010101010110001101010101;
		correct = 32'b00110010001110011100001010011101;
		#400 //-980127240000000.0 * -1.1031902e-23 = 1.0812667e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000011000100000011110000000110;
		b = 32'b10111001110010101010111100010001;
		correct = 32'b10111101011001000110001111111111;
		#400 //144.23447 * -0.00038658877 = -0.055759426
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100010111010110011100100110001;
		b = 32'b10100101001100001000111011010011;
		correct = 32'b01001000101000100011101010001101;
		#400 //-2.169553e+21 * -1.5313957e-16 = 332244.4
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001010110011011110001001001011;
		b = 32'b00111111100100011011110111000111;
		correct = 32'b11001010111010100110101110011001;
		#400 //-6746405.5 * 1.138604 = -7681484.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010000011011100000100100000011;
		b = 32'b01101110000001100011101100000100;
		correct = 32'b00111110111110011001111100101111;
		#400 //4.6944166e-29 * 1.0385584e+28 = 0.4875426
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011100011101111110000010110010;
		b = 32'b11010111011100010111010101000111;
		correct = 32'b00110100011010011100110000010110;
		#400 //-8.2015856e-22 * -265486000000000.0 = 2.1774062e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001100001011100111011110111101;
		b = 32'b01000010011001001111011111111100;
		correct = 32'b01001111000111000000101110100110;
		#400 //45735668.0 * 57.242172 = 2618009000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010001001000010000011001101100;
		b = 32'b00100001101000001010000010001100;
		correct = 32'b10110011010010100001000111111111;
		#400 //-43224842000.0 * 1.0884518e-18 = -4.7048157e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010010100000010000101110010101;
		b = 32'b01011011010001010001011110000110;
		correct = 32'b11101110010001101011001110001010;
		#400 //-277122550000.0 * 5.5476435e+16 = -1.537377e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110001101010001010011011011011;
		b = 32'b00010101111100111101111011011001;
		correct = 32'b11001000001000001010100100110010;
		#400 //-1.6702463e+30 * 9.849851e-26 = -164516.78
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000101001101001100001111000001;
		b = 32'b00011010001011111100000100001010;
		correct = 32'b00011111111110000011010000111111;
		#400 //2892.2346 * 3.6345088e-23 = 1.0511852e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110101000110101100000111001110;
		b = 32'b11011110110011000110001111000000;
		correct = 32'b01010100011101110001110101111010;
		#400 //-5.7651494e-07 * -7.363913e+18 = 4245405800000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111101100001101001111111100;
		b = 32'b01101010001101011000011111000011;
		correct = 32'b01110010011110101100011101001111;
		#400 //90535.97 * 5.4864172e+25 = 4.967181e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100000110010111100001101100001;
		b = 32'b10000000100001010000111011000101;
		correct = 32'b10100001110100111101000010000110;
		#400 //1.1746149e+20 * -1.2219419e-38 = -1.4353112e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010110111110110011100001110110;
		b = 32'b01010000000010011111111110001000;
		correct = 32'b11100111100001110110101111111010;
		#400 //-138109960000000.0 * 9260900000.0 = -1.2790226e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111101011011100100111001010000;
		b = 32'b11111010010010110100001101110111;
		correct = 32'b11111000001111010011011011100111;
		#400 //0.058180153 * -2.6385115e+35 = -1.5350901e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000011001001101001011101001;
		b = 32'b11010111111000001010110011011011;
		correct = 32'b01001000110010001101001100001101;
		#400 //-8.324564e-10 * -494066030000000.0 = 411288.4
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101101100011000110101111100011;
		b = 32'b01101111111110001111000110110110;
		correct = 32'b11011110000010001000110100011001;
		#400 //-1.5964069e-11 * 1.5408899e+29 = -2.459887e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011111111111001001101000110100;
		b = 32'b10001101100011101001001101110011;
		correct = 32'b10101110000011001010111100000111;
		#400 //3.6403836e+19 * -8.786923e-31 = -3.198777e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001010010000010001101001000001;
		b = 32'b01011111011111011110111000110000;
		correct = 32'b01101010001111111000101010011101;
		#400 //3163792.2 * 1.8297615e+19 = 5.7889854e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101111110010111100100001001111;
		b = 32'b01110011010100110001000110001010;
		correct = 32'b11100011101010000000010000001111;
		#400 //-3.7067813e-10 * 1.672257e+31 = -6.198691e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011111000010011010010110010;
		b = 32'b01100001001001010110010001000010;
		correct = 32'b11101101100100010111111100101001;
		#400 //-29518180.0 * 1.9068357e+20 = -5.6286317e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001110100011101000101110011000;
		b = 32'b01110000010101101110000111010000;
		correct = 32'b00111111011011110100110011011011;
		#400 //3.5140127e-30 * 2.6601113e+29 = 0.9347665
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111100100101011101101010011101;
		b = 32'b11010110011100011111011011101011;
		correct = 32'b01010011100011011010001101010111;
		#400 //-0.01829272 * -66510700000000.0 = 1216661600000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100001101000110110000100010;
		b = 32'b11010111110011011010000101000001;
		correct = 32'b11011100100100001110110000111101;
		#400 //721.6896 * -452184930000000.0 = -3.2633715e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010000110011000001011101001000;
		b = 32'b01111000110000000011011000101001;
		correct = 32'b11001010000110010011110010100100;
		#400 //-8.049968e-29 * 3.118811e+34 = -2510633.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111101000010100010111000101011;
		b = 32'b10101000010001110110000001011000;
		correct = 32'b01100101110101110011101111001000;
		#400 //-1.1479574e+37 * -1.106761e-14 = 1.27051445e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010011101100001001101100101011;
		b = 32'b00110101100111010011000111111110;
		correct = 32'b00001001110110001110001101001101;
		#400 //4.4581654e-27 * 1.1711961e-06 = 5.221386e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110011001101111000001001001110;
		b = 32'b10011101101000000101100110111110;
		correct = 32'b10010001011001011110001110001010;
		#400 //4.272652e-08 * -4.244444e-21 = -1.8135031e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000110110111101111001100000000;
		b = 32'b10100101000011101011111010111111;
		correct = 32'b00101100011110001010000111010001;
		#400 //-28537.5 * -1.2381164e-16 = 3.5332746e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011001100101100110010010000011;
		b = 32'b11000100101001110011010010010011;
		correct = 32'b00011110110001000111010011101000;
		#400 //-1.5550233e-23 * -1337.643 = 2.0800658e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111000010001010100100110001010;
		b = 32'b00110101000110100011100010101111;
		correct = 32'b10101101111011011011001111011000;
		#400 //-4.703695e-05 * 5.7451956e-07 = -2.7023647e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101011000110010010001011000001;
		b = 32'b01101011111101010101001111101011;
		correct = 32'b01010111100100101100000001110110;
		#400 //5.440475e-13 * 5.9316623e+26 = 322710620000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110101011111011001111000110110;
		b = 32'b10011100110000110000101101000111;
		correct = 32'b10010010110000010011101010101111;
		#400 //9.448007e-07 * -1.2906933e-21 = -1.2194479e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101001011010100011001010010101;
		b = 32'b00110110101000000111100101001001;
		correct = 32'b01100000100100101100111010010010;
		#400 //1.7695469e+25 * 4.782491e-06 = 8.4628425e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101011001000001100011100111111;
		b = 32'b11000010000001111100010111100001;
		correct = 32'b10101101101010101000101010110010;
		#400 //5.711993e-13 * -33.94324 = -1.9388356e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011101111000001101011001101100;
		b = 32'b10110001011001101111101010001011;
		correct = 32'b11001111110010101101110010110001;
		#400 //2.025157e+18 * -3.3611822e-09 = -6806921700.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110100110110011101100101100011;
		b = 32'b01011001000001001111111010011010;
		correct = 32'b01001110011000100101100110000000;
		#400 //4.057757e-07 * 2339664600000000.0 = 949379100.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000101001000110100101001101111;
		b = 32'b01101101110101101011110110110111;
		correct = 32'b10110011100010001111100100111011;
		#400 //-7.6778945e-36 * 8.307393e+27 = -6.378328e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010011111010011010110001001011;
		b = 32'b01000000011110110111111001111111;
		correct = 32'b01010100111001011000111101100100;
		#400 //2007236000000.0 * 3.9295957 = 7887625700000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111110001100110100111110001;
		b = 32'b10100110111000001010001001110000;
		correct = 32'b00011111001011100001101010011001;
		#400 //-2.3652772e-05 * -1.5587151e-15 = 3.6867934e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111011100101111010000001100101;
		b = 32'b11101001101001110101000001101111;
		correct = 32'b01100101110001100011001010001100;
		#400 //-0.004627275 * -2.5283806e+25 = 1.1699512e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000101001000100011100110001110;
		b = 32'b10011101111110010100001110010100;
		correct = 32'b00100011100111011111010011001110;
		#400 //-2595.5972 * -6.5979625e-21 = 1.7125653e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001010001000111101011101110110;
		b = 32'b00111110101001101110101110010000;
		correct = 32'b10001001010101011010100011110011;
		#400 //-7.888688e-33 * 0.32601595 = -2.5718382e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110111110000010011000110111;
		b = 32'b11011000001001000010000110110111;
		correct = 32'b01001111100111110001100100101010;
		#400 //-7.3954247e-06 * -721858840000000.0 = 5338453000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011101001111111111110110100110;
		b = 32'b11000010011010001000000000101010;
		correct = 32'b11100000001011100101110111111101;
		#400 //8.6464976e+17 * -58.12516 = -5.0257907e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001100001000101101000100000011;
		b = 32'b11001101001000110010001100010011;
		correct = 32'b11011001110011111000001011000111;
		#400 //42681356.0 * -171061550.0 = -7301139000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011110101001101000010011010011;
		b = 32'b10101100100010010010000101001101;
		correct = 32'b11001011101100100110010101111100;
		#400 //5.9994737e+18 * -3.8974713e-12 = -23382776.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111101000011111001010010010000;
		b = 32'b01011111011110100101010101111010;
		correct = 32'b11011101000011000110011100000101;
		#400 //-0.03505379 * 1.8038458e+19 = -6.323163e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010100111110110001110000100110;
		b = 32'b01100011000101111101000111011111;
		correct = 32'b11111000100101001110101101110111;
		#400 //-8628072300000.0 * 2.8005812e+21 = -2.4163617e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110010110001100110100100010000;
		b = 32'b10010111010110100100111111110001;
		correct = 32'b10001010101010010011001101101101;
		#400 //2.309801e-08 * -7.05405e-25 = -1.6293452e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011000101100110011111011110001;
		b = 32'b01100001010101011010001111111110;
		correct = 32'b01111010100101011001011000110001;
		#400 //1576663300000000.0 * 2.4631084e+20 = 3.8834924e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010101001011001100001110101100;
		b = 32'b10001110000111111110000110110110;
		correct = 32'b10100011110101111100101110110101;
		#400 //11872275000000.0 * -1.9706939e-30 = -2.339662e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100000101001101000111111001101;
		b = 32'b01011110111111101110000110100110;
		correct = 32'b01000000001001011101010101111110;
		#400 //2.8216653e-19 * 9.1830716e+18 = 2.5911555
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010000001110110100011101110111;
		b = 32'b10001100000010111011101001111000;
		correct = 32'b00011100110011000111000001101111;
		#400 //-12568092000.0 * -1.0764284e-31 = 1.3528651e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111000000001110001011000110111;
		b = 32'b11001000001111001001110100100000;
		correct = 32'b11000000110001110000111001110100;
		#400 //3.2207197e-05 * -193140.5 = -6.2205143
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010111101111100001001111000000;
		b = 32'b11100011111110100110110101101111;
		correct = 32'b11111100001110011111000010001010;
		#400 //417984070000000.0 * -9.239143e+21 = -3.8618145e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100010110001000100001100110101;
		b = 32'b00001101011011000100101000011101;
		correct = 32'b10110000101101010010011011000111;
		#400 //-1.8102023e+21 * 7.2812325e-31 = -1.3180504e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111000110010001111000010011;
		b = 32'b10000000110111110000010110001101;
		correct = 32'b10001000100001010110010010000100;
		#400 //39198.074 * -2.0481307e-38 = -8.028277e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000000010001110101001011100001;
		b = 32'b11001101100110001110110110111001;
		correct = 32'b10001110001010100110110111000011;
		#400 //6.550052e-39 * -320714530.0 = -2.1006966e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100110100100001011011001101001;
		b = 32'b01010100110100001001100110111001;
		correct = 32'b00111011111010111101011000110110;
		#400 //1.004145e-15 * 7167458000000.0 = 0.007197167
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010010101100000100110110010;
		b = 32'b10100101101111110111001111101011;
		correct = 32'b00100000101000000001001000100111;
		#400 //-0.0008164897 * -3.3211767e-16 = 2.7117067e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000101000011010011100001101010;
		b = 32'b01011010110100010101010101011100;
		correct = 32'b10100000011001101111010001001010;
		#400 //-6.64015e-36 * 2.9461062e+16 = -1.9562586e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111110111010011000001011010110;
		b = 32'b10000111000011011111111011010111;
		correct = 32'b00000110100000011000010110000100;
		#400 //-0.45607632 * -1.0682552e-34 = 4.872059e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111010100000110001010111000;
		b = 32'b00111100000100000100100011111101;
		correct = 32'b10110011111010101110010111100010;
		#400 //-1.2420751e-05 * 0.008806464 = -1.09382896e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010010101011000000110111000000;
		b = 32'b10100111010101101100101111101110;
		correct = 32'b10111010100100000101110010001101;
		#400 //369482530000.0 * -2.9809016e-15 = -0.001101391
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101010011000100101010111000111;
		b = 32'b10001011101000010100011110010010;
		correct = 32'b00110110100011101001011100111001;
		#400 //-6.8405577e+25 * -6.212263e-32 = 4.2495344e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000010011010001100001101010110;
		b = 32'b01100001001010010100100000000100;
		correct = 32'b11100100000110011110101001101110;
		#400 //-58.190758 * 1.9516806e+20 = -1.1356977e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000001111101010000101010000011;
		b = 32'b10000011100011000001001010111100;
		correct = 32'b10000110000001100001001110101110;
		#400 //30.630133 * -8.232762e-37 = -2.5217057e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111101101000110101001010001100;
		b = 32'b01111111010100101111110110011101;
		correct = 32'b11111101100001101001101110000100;
		#400 //-0.07974729 * 2.8045471e+38 = -2.2365504e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101001000011110001110000011100;
		b = 32'b10100001111001101100001110101110;
		correct = 32'b11001011100000010000000010100101;
		#400 //1.0813071e+25 * -1.5637202e-18 = -16908618.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001100111010110110011001010111;
		b = 32'b10011001101110001000001111101110;
		correct = 32'b10100111001010011010101011011111;
		#400 //123417270.0 * -1.907844e-23 = -2.354609e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100101110110011110100010001110;
		b = 32'b10110010011111101111001111011010;
		correct = 32'b01011000110110010000010001001110;
		#400 //-1.28630425e+23 * -1.4840191e-08 = 1908900100000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100110000110100011000000011110;
		b = 32'b01011011001110111101111000111101;
		correct = 32'b11000001111000100100111000000001;
		#400 //-5.3494694e-16 * 5.2880174e+16 = -28.288088
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110110111000000001010111100110;
		b = 32'b01000000000001101010001001100011;
		correct = 32'b00110111011010111011001100110110;
		#400 //6.6782695e-06 * 2.1036613 = 1.4048817e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000101010100011000100011110101;
		b = 32'b10001111000111101010101010100001;
		correct = 32'b10010101000000011101111000110000;
		#400 //3352.5598 * -7.822863e-30 = -2.6226618e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000000000000100111001111110101;
		b = 32'b00011001011010111111011111100000;
		correct = 32'b00011001111100000111110110000100;
		#400 //2.0383275 * 1.2199273e-23 = 2.4866114e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110011010001100010111010101100;
		b = 32'b00011100001101100000111111011111;
		correct = 32'b10010000000011001111000101111000;
		#400 //-4.6142915e-08 * 6.023926e-22 = -2.7796152e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001110000111011000111101001101;
		b = 32'b10011001000110100100000011000000;
		correct = 32'b00100111101111011110000000011101;
		#400 //-660853570.0 * -7.9746896e-24 = 5.270102e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100110101001000010111000001000;
		b = 32'b10100000001001011011101001000001;
		correct = 32'b11000111010101001001001000111101;
		#400 //3.876586e+23 * -1.403767e-19 = -54418.24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010110001110111000010000101111;
		b = 32'b01011110110011011100100110000011;
		correct = 32'b00110101100101101011110001110100;
		#400 //1.514745e-25 * 7.4142636e+18 = 1.1230718e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101111101010000101001111101011;
		b = 32'b01111110110111001100100101011001;
		correct = 32'b11101111000100010010110010000010;
		#400 //-3.061865e-10 * 1.4673781e+38 = -4.4929133e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100000111101110000010011110000;
		b = 32'b01011000100100001111001111110011;
		correct = 32'b01111010000010111101111000101011;
		#400 //1.4239692e+20 * 1275019400000000.0 = 1.8155884e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101000111100000111010011100111;
		b = 32'b11010111111001000100010101000100;
		correct = 32'b01000001010101100110100100101101;
		#400 //-2.6696051e-14 * -501972300000000.0 = 13.400678
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001101100101101101010001001010;
		b = 32'b00101100100011011001101100011010;
		correct = 32'b00111010101001101101110010011101;
		#400 //316311870.0 * 4.0246808e-12 = 0.0012730543
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000000011000011101101000101001;
		b = 32'b01111101010111000101001011100010;
		correct = 32'b01111110010000100110000010011010;
		#400 //3.5289404 * 1.8303782e+37 = 6.4592954e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100100100111011010000111101000;
		b = 32'b11010100000010110011100001100110;
		correct = 32'b01111001001010110111001101000110;
		#400 //-2.3262443e+22 * -2391786700000.0 = 5.56388e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001101111100011010010110111100;
		b = 32'b11000001100101100000100001011001;
		correct = 32'b00010000000011011001111011111101;
		#400 //-1.4892671e-30 * -18.754076 = 2.7929827e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010110011100010010100011111;
		b = 32'b10101010100100010001001011110010;
		correct = 32'b00100101111010011010010010010000;
		#400 //-0.0015727616 * -2.577032e-13 = 4.053057e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111001001010101110010100001111;
		b = 32'b00111000010100110011101110011001;
		correct = 32'b00110010000011010000001010010100;
		#400 //0.00016297794 * 5.0361825e-05 = 8.207866e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101100110000100000110110010000;
		b = 32'b10011101010111010110010011010001;
		correct = 32'b10001010101001111101001000100001;
		#400 //5.5153174e-12 * -2.9301227e-21 = -1.6160557e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101100001001011011000001011010;
		b = 32'b00010101000110011100111001100110;
		correct = 32'b01000001110001110001011111110111;
		#400 //8.012222e+26 * 3.1060924e-26 = 24.886702
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110110110011010101001110000111;
		b = 32'b00101010111101111111000101101000;
		correct = 32'b01100010010001101101110100110110;
		#400 //2.0822558e+33 * 4.4043523e-13 = 9.170988e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100011110111011111111011110100;
		b = 32'b00111100011011000011001111011011;
		correct = 32'b00100000110011001101010000000001;
		#400 //2.4068845e-17 * 0.01441666 = 3.4699237e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011000101001111110110110101101;
		b = 32'b11011110011011111100001100101000;
		correct = 32'b00110111100111010100011011101001;
		#400 //-4.340848e-24 * -4.3191741e+18 = 1.8748879e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100110000001111000011001001101;
		b = 32'b00011100010001001110100100011101;
		correct = 32'b00000010110100000111110001110111;
		#400 //4.7019545e-16 * 6.515225e-22 = 3.0634292e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011000011010001011110111010100;
		b = 32'b01001111100001110001111001011100;
		correct = 32'b00101000011101011010111101101001;
		#400 //3.0081136e-24 * 4533827600.0 = 1.3638268e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110010001011011001100111011110;
		b = 32'b00001110111101100011001011111111;
		correct = 32'b01000001101001101111010001110000;
		#400 //3.438523e+30 * 6.069279e-30 = 20.869354
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111101110001010101100110100101;
		b = 32'b10101000000001010000010010100001;
		correct = 32'b00100110010011010001011001001000;
		#400 //-0.09636239 * -7.383987e-15 = 7.115386e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110110010110001010101111000001;
		b = 32'b00000011010011101000001101101110;
		correct = 32'b10111010001011101100100101110010;
		#400 //-1.09865206e+33 * 6.0688833e-37 = -0.0006667591
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110001000010101011010100111101;
		b = 32'b00100110000000100011011011101111;
		correct = 32'b10010111100011010001101110011001;
		#400 //-2.0184665e-09 * 4.517726e-16 = -9.118878e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110100111110111110001000101110;
		b = 32'b10111010001110111111110101011111;
		correct = 32'b01101111101110001111011110000100;
		#400 //-1.5965014e+32 * -0.0007171239 = 1.1448894e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100110010101011101011100100;
		b = 32'b01000111101111000001001011111001;
		correct = 32'b01001101000101001111000001000110;
		#400 //1621.8403 * 96293.945 = 156173400.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010111110010000111011111110110;
		b = 32'b10000100001011001111110101000011;
		correct = 32'b00011100100001110111011011101100;
		#400 //-440835100000000.0 * -2.0334795e-36 = 8.964291e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001100001101100110111010010001;
		b = 32'b10101101011100000110101100110001;
		correct = 32'b10111010001010110101010000001011;
		#400 //47823428.0 * -1.3666222e-11 = -0.00065356557
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001100101011100011011000010000;
		b = 32'b01000111100011111001110101111000;
		correct = 32'b11010100110000110111011010111000;
		#400 //-91336830.0 * 73530.94 = -6716083000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101010001000100111010100101001;
		b = 32'b00100101110101010110001101000010;
		correct = 32'b01010000100001110110101001111000;
		#400 //4.9099814e+25 * 3.701687e-16 = 18175214000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101100110000100010011001100000;
		b = 32'b10100110001100111111101001001110;
		correct = 32'b01010011100010000111111010101010;
		#400 //-1.8777026e+27 * -6.2442327e-16 = 1172481200000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001111000011101110111011000111;
		b = 32'b11111111110001011101110000111001;
		correct = 32'b11111111110001011101110000111001;
		#400 //2398013200.0 * nan = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011111000111100010000001000110;
		b = 32'b11101111011010001110001011000010;
		correct = 32'b01001111000011111101100101010000;
		#400 //-3.3484497e-20 * -7.2074656e+28 = 2413383700.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010101001101111110111010010001;
		b = 32'b01011101111010010110101101100010;
		correct = 32'b10110011101001111011010101001001;
		#400 //-3.714475e-26 * 2.1024556e+18 = -7.809519e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011010010101000101100000100100;
		b = 32'b11010100111001110010001110110010;
		correct = 32'b11101111101111111011100100100100;
		#400 //1.4942402e+16 * -7941890500000.0 = -1.1867092e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100011010011111100110110110110;
		b = 32'b00010010110000001101011101011110;
		correct = 32'b00110110100111001000100100011011;
		#400 //3.833299e+21 * 1.2169996e-27 = 4.6651235e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110001010100000010100010001111;
		b = 32'b10011110010001011111100011110110;
		correct = 32'b10010000001000001111100110100101;
		#400 //3.0291039e-09 * -1.0480577e-20 = -3.1746755e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001001011110101011000100110100;
		b = 32'b01100010100100011110111000111101;
		correct = 32'b10101100100011101110011110101011;
		#400 //-3.0175976e-33 * 1.3459724e+21 = -4.061603e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010110001010111001010110010111;
		b = 32'b10000000010001101110000101000011;
		correct = 32'b00010110101111100000011110001011;
		#400 //-47164743000000.0 * -6.509293e-39 = 3.0700916e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010001101111100000101011100111;
		b = 32'b00110111110111111111001101000100;
		correct = 32'b10001010001001100100000000010110;
		#400 //-2.9983433e-28 * 2.6696951e-05 = -8.0046625e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011111001111000111110000100100;
		b = 32'b01010000000001010100101010110100;
		correct = 32'b10101111110001000100011011111110;
		#400 //-3.9913235e-20 * 8945062000.0 = -3.5702635e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000100011000111011100001001101;
		b = 32'b00110111010000110010011111001001;
		correct = 32'b10111100001011011001100011000111;
		#400 //-910.8797 * 1.1632169e-05 = -0.010595507
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011011101101101100111010111000;
		b = 32'b10111100001100110001011101000100;
		correct = 32'b00011000011111111100011001010000;
		#400 //-3.0242963e-22 * -0.01093084 = 3.30581e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000101011101110100100100100000;
		b = 32'b01101000011101000000010001100101;
		correct = 32'b10101110011010111011010111110001;
		#400 //-1.1627315e-35 * 4.609354e+24 = -5.359441e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101001111000100101110101001000;
		b = 32'b01000010101101100001101011000110;
		correct = 32'b11101101001000010000010111111110;
		#400 //-3.4207218e+25 * 91.05229 = -3.1146457e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100101101001011100111010001101;
		b = 32'b10110110101001011001010100011001;
		correct = 32'b11011100110101100111110101100101;
		#400 //9.787508e+22 * -4.9347404e-06 = -4.8298814e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001100100110010010101100100000;
		b = 32'b10001011001010110000001110000101;
		correct = 32'b00011000010011001010001111010011;
		#400 //-80304380.0 * -3.293605e-32 = 2.6449092e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101110100111011010000000101100;
		b = 32'b10101101101010101010110100010100;
		correct = 32'b00011100110100100010110111011110;
		#400 //-7.1679856e-11 * -1.9403625e-11 = 1.3908491e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010011110100010000101110010011;
		b = 32'b11001110100100101000101110100110;
		correct = 32'b01100010111011110101010101000101;
		#400 //-1795684700000.0 * -1229312800.0 = 2.2074581e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111101010110010001011111001111;
		b = 32'b10100111101111011010101000101101;
		correct = 32'b00100101101000001101011011100100;
		#400 //-0.05300122 * -5.2642543e-15 = 2.790119e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010111101110001101001000100100;
		b = 32'b11011110010111001110000101011010;
		correct = 32'b00110110100111110111011101001001;
		#400 //-1.1943768e-24 * -3.9790254e+18 = 4.752456e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100110000111000100011001101010;
		b = 32'b00000011110110100000011010101110;
		correct = 32'b10101010100001010001100000001010;
		#400 //-1.8449702e+23 * 1.2814422e-36 = -2.3642226e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110000100100111100100111011100;
		b = 32'b11000001001110001011110110011000;
		correct = 32'b10110010010101010100110100010100;
		#400 //1.075303e-09 * -11.546288 = -1.2415757e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100101101100110111011110011110;
		b = 32'b10101010101100101001011101111111;
		correct = 32'b11010000111110100110011011000001;
		#400 //1.0593877e+23 * -3.1724273e-13 = -33608305000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010011010001101011010101010100;
		b = 32'b10111011010111110011110000001011;
		correct = 32'b01001111001011010100011010001111;
		#400 //-853445700000.0 * -0.0034062888 = 2907082500.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001111000111111111000000000001;
		b = 32'b01001100101001100101001011111101;
		correct = 32'b10011100010011111101001011110011;
		#400 //-7.885528e-30 * 87201770.0 = -6.87632e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110100110001000100100111001101;
		b = 32'b00100111111001111111110100101010;
		correct = 32'b10011101001100011110000010110101;
		#400 //-3.6561542e-07 * 6.438986e-15 = -2.3541926e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010110011101000100000001001011;
		b = 32'b00010111111111111111010101001000;
		correct = 32'b10101110111101000011011000010001;
		#400 //-67139243000000.0 * 1.6540906e-24 = -1.11054395e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101100101101011101101000100010;
		b = 32'b00100101010010010000011110010001;
		correct = 32'b10010010100011101100110110100101;
		#400 //-5.168547e-12 * 1.7436535e-16 = -9.012155e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011101110001100010110010000100;
		b = 32'b10101111100000001111000110100001;
		correct = 32'b10001101110001111010001010011101;
		#400 //5.245619e-21 * -2.3454752e-10 = -1.230347e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010010010000110001011011110000;
		b = 32'b10101111110010110010111011001011;
		correct = 32'b11000010100110101101011011011001;
		#400 //209475860000.0 * -3.6958733e-10 = -77.419624
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011111000101110001100011000000;
		b = 32'b10110010111010111100110111101011;
		correct = 32'b11010010100010110010110101000010;
		#400 //1.0887663e+19 * -2.7451241e-08 = -298879880000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001111010010111011010011100001;
		b = 32'b01000000110100000111101111100010;
		correct = 32'b01010000101001011110010110001011;
		#400 //3417629000.0 * 6.5151224 = 22266272000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101100001001000011101100101010;
		b = 32'b00110110011100100001100011110011;
		correct = 32'b11100011000110110100111111101111;
		#400 //-7.941729e+26 * 3.6075332e-06 = -2.8650052e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100100110100101100111011111000;
		b = 32'b01111111011001011111001001010011;
		correct = 32'b01100100101111010101101010110000;
		#400 //9.14236e-17 * 3.0565143e+38 = 2.7943755e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000011110111001001100011111001;
		b = 32'b00101010001000001110000011011000;
		correct = 32'b00101110100010101010000101011100;
		#400 //441.1951 * 1.4288863e-13 = 6.3041766e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110011000011000111100000001101;
		b = 32'b11000010001100101111010010010001;
		correct = 32'b10110101110001000110001101010110;
		#400 //3.2705476e-08 * -44.738834 = -1.4632049e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001010111101011000101010011110;
		b = 32'b10110001011101001000100110010110;
		correct = 32'b10111100111010101000110000010110;
		#400 //8045903.0 * -3.5584882e-09 = -0.028631251
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000110011111111111100001000001;
		b = 32'b10110011111000000100100100000101;
		correct = 32'b10111010111000000100001000111100;
		#400 //16382.063 * -1.0444095e-07 = -0.0017109583
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001011000001111010011011011101;
		b = 32'b10111101010000011101101110011010;
		correct = 32'b11001000110011010111001001010100;
		#400 //8890077.0 * -0.04732857 = -420754.62
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100111100101001111010110011100;
		b = 32'b01001010010110000111110110011000;
		correct = 32'b01110010011110111111000010100000;
		#400 //1.4068819e+24 * 3546982.0 = 4.9901847e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100000101010011011011101100010;
		b = 32'b01101100110101100001110000000111;
		correct = 32'b11001110000011011111000111100001;
		#400 //-2.8751066e-19 * 2.0707398e+27 = -595359800.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000001110001110111011011000010;
		b = 32'b11110000011011001001001101011010;
		correct = 32'b00110010101110000101010001001010;
		#400 //-7.3271464e-38 * -2.928664e+29 = 2.145875e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111011011000000001011001000100;
		b = 32'b10001101100011101001011111100111;
		correct = 32'b00001001011110011010001010100010;
		#400 //-0.003419296 * -8.787995e-31 = 3.0048754e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010101010011000101100110110100;
		b = 32'b00110111010000100101000101101111;
		correct = 32'b00001101000110110001110011111011;
		#400 //4.1268235e-26 * 1.1582261e-05 = 4.7797947e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011111110001011011111001011100;
		b = 32'b10101100110010001000110111101010;
		correct = 32'b00001101000110101110101001010110;
		#400 //-8.374767e-20 * -5.7000975e-12 = 4.7736985e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000101111110011100110000100110;
		b = 32'b11011111011011111110101101110111;
		correct = 32'b10100101111010100001101101011010;
		#400 //2.349084e-35 * -1.7288042e+19 = -4.0611063e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101101011100010111101001001100;
		b = 32'b01011101110100011101011101000000;
		correct = 32'b01001011110001011110111111100010;
		#400 //1.3726419e-11 * 1.8900781e+18 = 25944004.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001001011001010110100011001111;
		b = 32'b10000000010001100101110111111101;
		correct = 32'b10001001111111000011101110001010;
		#400 //939660.94 * -6.462201e-39 = -6.0722784e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000111001110001111010101110011;
		b = 32'b11100111101011000110111111110011;
		correct = 32'b01101111011110010010101110010111;
		#400 //-47349.45 * -1.6286243e+24 = 7.7114464e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111001111110111011010000010111;
		b = 32'b00100111101001100100101010101000;
		correct = 32'b00100010001000111000000000101110;
		#400 //0.00048008628 * 4.61552e-15 = 2.2158477e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101010011101101011001111010100;
		b = 32'b01111100101001110010010111100001;
		correct = 32'b01100111101000010001001111010000;
		#400 //2.191158e-13 * 6.943055e+36 = 1.521333e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000011000001011111001011110010;
		b = 32'b10100101100011110101100000100011;
		correct = 32'b00101001000101100000000110100110;
		#400 //-133.949 * -2.486627e-16 = 3.330812e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101111110011111110000011101110;
		b = 32'b01000101011010110010000111100100;
		correct = 32'b00110101101111101110111100000000;
		#400 //3.7812903e-10 * 3762.1182 = 1.4225661e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101100011101101111010010001011;
		b = 32'b00100011011111111011000010100011;
		correct = 32'b00010000011101101010011111111100;
		#400 //3.5094451e-12 * 1.3860982e-17 = 4.8644356e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100001111111000010101011110111;
		b = 32'b00111100101001011011001111010100;
		correct = 32'b11011111001000110011100011010100;
		#400 //-5.8145943e+20 * 0.02022735 = -1.1761384e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001110010000110001111011001000;
		b = 32'b01010001011001110001110010101000;
		correct = 32'b11100000001100000010011010011110;
		#400 //-818393600.0 * 62038640000.0 = -5.0772025e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000001001010110100010110011;
		b = 32'b01000111101000001101011111110101;
		correct = 32'b10111000010011111101100111110010;
		#400 //-6.0175437e-10 * 82351.914 = -4.9555623e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111100101110111010011111000110;
		b = 32'b01111101100000011001101001100011;
		correct = 32'b01111010101111100000000101101101;
		#400 //0.022907149 * 2.1534004e+37 = 4.9328266e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011000101010100001001000101100;
		b = 32'b10111010001100100110011011111111;
		correct = 32'b10010011011011010000101000011110;
		#400 //4.396232e-24 * -0.0006805509 = -2.9918594e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001011101101100011110111010011;
		b = 32'b01001100011110100110101101110011;
		correct = 32'b10011000101100100100010011011110;
		#400 //-7.019687e-32 * 65646028.0 = -4.608146e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010111011100011100001111101110;
		b = 32'b01010100101011011110100011011011;
		correct = 32'b01101100101001000011110101010000;
		#400 //265823810000000.0 * 5975488000000.0 = 1.588427e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101101100000011010110110110100;
		b = 32'b10001100111110010011000111111111;
		correct = 32'b00111010111111000111011010001111;
		#400 //-5.016695e+27 * -3.8394615e-31 = 0.0019261407
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010011000000101011110000111001;
		b = 32'b00011110101011101011101010111011;
		correct = 32'b10110010001100100111011010010110;
		#400 //-561503600000.0 * 1.8500197e-20 = -1.0387927e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000111101101110001110011011110;
		b = 32'b11000100001001000010010011101101;
		correct = 32'b10001100011010101101000111010000;
		#400 //2.7551746e-34 * -656.57697 = -1.8089842e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011100011000001001110000001;
		b = 32'b00100001011000111010110010101100;
		correct = 32'b10101101011110010010011110001101;
		#400 //-18360066.0 * 7.713912e-19 = -1.4162793e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001010011101011001000010100000;
		b = 32'b11011100011110101101100110110000;
		correct = 32'b10100111011100001010000000001101;
		#400 //1.1823522e-32 * -2.8243238e+17 = -3.3393454e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111001011110011001000110111010;
		b = 32'b11010101100111110011100101001001;
		correct = 32'b11001111100110110011100101011011;
		#400 //0.00023800778 * -21883548000000.0 = -5208454700.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000101100011000101110010100010;
		b = 32'b10101000111000111110001011101011;
		correct = 32'b10101110111110011110010100011101;
		#400 //4491.579 * -2.5300473e-14 = -1.1363908e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110011101100101001011111100111;
		b = 32'b11000111011110010001000111100110;
		correct = 32'b11111011101011011100001000111100;
		#400 //2.829925e+31 * -63761.9 = -1.8044138e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100001110010010101100101110100;
		b = 32'b00100010111111111110101101000011;
		correct = 32'b10000101010010010100100100100100;
		#400 //-1.3643968e-18 * 6.936698e-18 = -9.4644084e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000111111010000000101010110101;
		b = 32'b01011101001111010011010111001101;
		correct = 32'b10100101101010111000000010101100;
		#400 //-3.4913773e-34 * 8.521268e+17 = -2.9750963e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011000100111011101110111110110;
		b = 32'b10101010100010110001000010000011;
		correct = 32'b01000011101010111000001101100110;
		#400 //-1388613100000000.0 * -2.4702817e-13 = 343.02655
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110111010000010000000010001101;
		b = 32'b01000000110000010100000101001101;
		correct = 32'b00111000100100011011001010100101;
		#400 //1.1503825e-05 * 6.0392213 = 6.947414e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010010010101101010000010111011;
		b = 32'b00100100110110011001000100000000;
		correct = 32'b10110111101101100110011111010000;
		#400 //-230454900000.0 * 9.435439e-17 = -2.1744432e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011001100110001111010100111000;
		b = 32'b00101010101100010111011000011011;
		correct = 32'b01000100110101000001000000111010;
		#400 //5381727000000000.0 * 3.1523468e-13 = 1696.5071
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100010000001010000011101110110;
		b = 32'b01100000100010001001010000111001;
		correct = 32'b01000011000011011111000111111001;
		#400 //1.802881e-18 * 7.873243e+19 = 141.9452
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000010111111101001010101000110;
		b = 32'b11011011011000000110100001101101;
		correct = 32'b01011110110111110010101001110110;
		#400 //-127.29155 * -6.316521e+16 = 8.0403976e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100010001111010010000011110010;
		b = 32'b11001001100100100000100011011000;
		correct = 32'b11101100010101111100011010100101;
		#400 //8.7220215e+20 * -1196315.0 = -1.0434285e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101000111110011110001100110111;
		b = 32'b10110001000010011000001100010000;
		correct = 32'b00011010100001100011101010000111;
		#400 //-2.7743092e-14 * -2.0010624e-09 = 5.551566e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111101010000011101011001001100;
		b = 32'b10010010111101001010110111111111;
		correct = 32'b10010000101110010100001111111111;
		#400 //0.04732351 * -1.5441458e-27 = -7.30744e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011100111110100011000111000100;
		b = 32'b00000100100011110100100100011100;
		correct = 32'b00100010000011000000100101000000;
		#400 //5.633877e+17 * 3.368628e-36 = 1.8978435e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101111001011101101010100011110;
		b = 32'b10111111000110111101010111101010;
		correct = 32'b11101110110101001101101001000001;
		#400 //5.4108035e+28 * -0.6087328 = -3.2937337e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111101011100110101010110100010;
		b = 32'b10110111110101101011001111011111;
		correct = 32'b01110101110011000001010010001110;
		#400 //-2.021544e+37 * -2.5594547e-05 = 5.17405e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101100000000010001101111011110;
		b = 32'b10101100111000110100100011010001;
		correct = 32'b10011001011001010100000011011110;
		#400 //1.8347472e-12 * -6.4598123e-12 = -1.1852122e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011000100011100010010101101111;
		b = 32'b10001000110011011011111011010101;
		correct = 32'b00100001111001000111101111100000;
		#400 //-1250331400000000.0 * -1.2382853e-33 = 1.548267e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001001011100000000100001100000;
		b = 32'b01010011100001000010001111011000;
		correct = 32'b11011101011101111100101111011010;
		#400 //-983174.0 * 1135074100000.0 = -1.1159753e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101000001011110011001100101111;
		b = 32'b01110010101011001101100000010100;
		correct = 32'b01011011011011001001010010001001;
		#400 //9.72555e-15 * 6.8470584e+30 = 6.659141e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010011110111010010000111011110;
		b = 32'b11000001001101001101111010011010;
		correct = 32'b00010101100111000011110000011000;
		#400 //-5.582164e-27 * -11.304346 = 6.310271e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000111110010011010000101010100;
		b = 32'b11000011000111011111110001111010;
		correct = 32'b10001011011110001101110110010111;
		#400 //3.0337939e-34 * -157.98624 = -4.7929768e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111000010010000001011011100001;
		b = 32'b11111001101110111101111111001111;
		correct = 32'b01110010100100101101011110100100;
		#400 //-4.7705023e-05 * -1.2193736e+35 = 5.8170246e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100111100101100011110100100011;
		b = 32'b10110001000011110011011111011101;
		correct = 32'b00011001001010000001100111011111;
		#400 //-4.169965e-15 * -2.0840993e-09 = 8.690621e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010110001011101001010010101011;
		b = 32'b11001011101000110011110100101001;
		correct = 32'b10100010010111101010010010111101;
		#400 //1.410252e-25 * -21396050.0 = -3.0173822e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000101110001111111011001001;
		b = 32'b11110010000100101110101100010000;
		correct = 32'b01100011010101000101011001011000;
		#400 //-1.3460176e-09 * -2.910015e+30 = 3.9169315e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110111111101100101101011110000;
		b = 32'b00011110100000011001001111100110;
		correct = 32'b11010110111110010110010001001101;
		#400 //-9.993355e+33 * 1.3719576e-20 = -137104590000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101000010010110000110000010000;
		b = 32'b01000000101110100110100011110000;
		correct = 32'b00101001100100111101100111111111;
		#400 //1.1271379e-14 * 5.8253098 = 6.565928e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001100100101010001010000011110;
		b = 32'b01101110001010110100000111010000;
		correct = 32'b11111011010001110111010110000111;
		#400 //-78160110.0 * 1.3250375e+28 = -1.0356508e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110100011001011001001101010111;
		b = 32'b10010101001111111100001100001011;
		correct = 32'b00001010001010111111011111010111;
		#400 //-2.1380889e-07 * -3.8726005e-26 = 8.279964e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101110011011101010100010101000;
		b = 32'b10100100001000001011110010101111;
		correct = 32'b10010011000101011101100101010000;
		#400 //5.426473e-11 * -3.485429e-17 = -1.8913587e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001110101111001011111001111011;
		b = 32'b01001111000001101110011100110000;
		correct = 32'b00011110010001101110110001001111;
		#400 //4.6529004e-30 * 2263298000.0 = 1.05309e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111100101100011101010010100010;
		b = 32'b10100000110010011110110110110010;
		correct = 32'b01011110000011000100010100010001;
		#400 //-7.386794e+36 * -3.4208018e-19 = 2.526876e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010001011111111101100011001010;
		b = 32'b01011010101101000110010111001101;
		correct = 32'b11101100101101000100101000101011;
		#400 //-68678360000.0 * 2.5388713e+16 = -1.7436552e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000101000011101100011111011010;
		b = 32'b01001000101111111100000110111110;
		correct = 32'b11001110010101011110011001010101;
		#400 //-2284.4907 * 392717.94 = -897160500.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010101011001100100000111000010;
		b = 32'b01111111111101001100010001111100;
		correct = 32'b01111111111101001100010001111100;
		#400 //15823131000000.0 * nan = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110010011000001110011011000101;
		b = 32'b11000100110011011101110010110011;
		correct = 32'b10110111101101001101101010101111;
		#400 //1.3090987e-08 * -1646.8969 = -2.1559505e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110100111001101001001000110100;
		b = 32'b01001010111101011111110001100001;
		correct = 32'b01000000010111011000110100111011;
		#400 //4.2947215e-07 * 8060464.5 = 3.461745
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000110010110001111100011001101;
		b = 32'b01110010000100101010010110011110;
		correct = 32'b00111000111110001001010010000110;
		#400 //4.0807875e-35 * 2.904642e+30 = 0.00011853226
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100101101000100100001110100100;
		b = 32'b00101110011001100000110010110111;
		correct = 32'b01010100100100011101000011010101;
		#400 //9.578389e+22 * 5.230724e-11 = 5010191000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001010100111011100001011111010;
		b = 32'b01011101010001101000001000100111;
		correct = 32'b01101000011101001010101000000101;
		#400 //5169533.0 * 8.940024e+17 = 4.621575e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110110000111101110101011101010;
		b = 32'b10011101010010111000110110000101;
		correct = 32'b10010011111111001011100001000011;
		#400 //2.3680573e-06 * -2.693999e-21 = -6.379544e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111011110111110001101111011100;
		b = 32'b00001011011000000010101011011001;
		correct = 32'b10000111110000110101110110111000;
		#400 //-0.006808741 * 4.3173066e-32 = -2.9395422e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110011101000100001000011101;
		b = 32'b00001000111001010011110111100011;
		correct = 32'b00000111110110101011101000110000;
		#400 //0.23853345 * 1.3796986e-33 = 3.2910426e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001011111110010101011101001111;
		b = 32'b00010000000101111010110111010011;
		correct = 32'b00011100100100111011101111001101;
		#400 //32681630.0 * 2.9913408e-29 = 9.776189e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001111010100001110110010000010;
		b = 32'b01110010111001110110010100000101;
		correct = 32'b01000010101111001101011111011011;
		#400 //1.03007415e-29 * 9.166485e+30 = 94.42159
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110100001100011011101001100111;
		b = 32'b00101111111101001101010100010110;
		correct = 32'b10100100101010011111100110011010;
		#400 //-1.6552222e-07 * 4.4534748e-10 = -7.371491e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100111001100000001111101110110;
		b = 32'b11001101101100100010101011001101;
		correct = 32'b11110101011101010010011010100100;
		#400 //8.3171685e+23 * -373643680.0 = -3.1076574e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001011001111001000011111100001;
		b = 32'b11011001010001100011111110101100;
		correct = 32'b10100101000100011111111111111100;
		#400 //3.6309707e-32 * -3487628300000000.0 = -1.2663476e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001111110000000011111001110110;
		b = 32'b01101000110111110010000100000110;
		correct = 32'b11111001001001111000111100110101;
		#400 //-6450638000.0 * 8.429575e+24 = -5.4376135e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001110000100110011011101101100;
		b = 32'b01010100111101111011010100100110;
		correct = 32'b01100011100011100111001010100101;
		#400 //617470700.0 * 8511168700000.0 = 5.2553973e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001011110111001100011000101100;
		b = 32'b11001111110101001100100010011011;
		correct = 32'b10011100001101111000000100011101;
		#400 //8.5039093e-32 * -7139833300.0 = -6.0716496e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011011100000011111001000001001;
		b = 32'b11011110000100111110010001100110;
		correct = 32'b11111010000101100010001111010101;
		#400 //7.3152785e+16 * -2.6641887e+18 = -1.9489282e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111101111110001100010111100000;
		b = 32'b00100010001110111001000100111010;
		correct = 32'b10100000101101100100010110101011;
		#400 //-0.12147117 * 2.5420108e-18 = -3.0878102e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101101101001000000000010001011;
		b = 32'b11000010110111101010111110111110;
		correct = 32'b11110001000011101010100100001111;
		#400 //6.344525e+27 * -111.34325 = -7.0642e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110010011010110101011011001110;
		b = 32'b10010011000000101011011000111100;
		correct = 32'b11000101111100000101001100110111;
		#400 //4.6613707e+30 * -1.6498155e-27 = -7690.402
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010111101111110010001000010110;
		b = 32'b00111010010000111000001000111000;
		correct = 32'b00010010100100011111100000110000;
		#400 //1.235169e-24 * 0.0007458064 = 9.211969e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100010011110011000101011111001;
		b = 32'b01101100010110110100101011000011;
		correct = 32'b11001111010101011100001011000011;
		#400 //-3.3819364e-18 * 1.0604312e+27 = -3586311000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011100111011110110100011011110;
		b = 32'b01011011111010100111101011000011;
		correct = 32'b00111001010110110100100010101001;
		#400 //1.5842801e-21 * 1.32000245e+17 = 0.00020912536
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011011011010001010110111000101;
		b = 32'b01111010001101100101010011011000;
		correct = 32'b11010110001001011011100010100111;
		#400 //-1.9246738e-22 * 2.3667972e+35 = -45553124000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000010000110011100100011001010;
		b = 32'b00110111001100011101010000100001;
		correct = 32'b10111001110101011010011010000100;
		#400 //-38.446083 * 1.0599412e-05 = -0.0004075059
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010001110100000011001111010110;
		b = 32'b00001101100001010110100010100010;
		correct = 32'b10011111110110010000000000001110;
		#400 //-111777860000.0 * 8.221947e-31 = -9.1903165e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111100110100100011100011101110;
		b = 32'b00111001001001101010110001110000;
		correct = 32'b00110110100010001101111010000101;
		#400 //0.025661912 * 0.00015895232 = 4.0790205e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001110011000100000110001011011;
		b = 32'b01011101100000110100000010010001;
		correct = 32'b01101100011001111100101010101011;
		#400 //948115140.0 * 1.1822148e+18 = 1.12087575e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111101110001001101011100110100;
		b = 32'b11100010101101101100101101001010;
		correct = 32'b01100001000011001000110101001111;
		#400 //-0.09611359 * -1.685978e+21 = 1.620454e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111111000100110101100100011111;
		b = 32'b00110000110101000011010000101111;
		correct = 32'b00110000011101000100011110101110;
		#400 //0.57557863 * 1.5439862e-09 = 8.8868546e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101010111001000111011001010111;
		b = 32'b11000101010011011000101010110000;
		correct = 32'b11110000101101110110111010001001;
		#400 //1.3809697e+26 * -3288.668 = -4.541551e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100001111101110000111110100001;
		b = 32'b11100111101011010110101011100011;
		correct = 32'b01001010001001110101110010110111;
		#400 //-1.6741508e-18 * -1.6378822e+24 = 2742061.8
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010001101000011001001001101010;
		b = 32'b11011001011010100001110000100001;
		correct = 32'b11101011100100111100000110010110;
		#400 //86743270000.0 * -4118504500000000.0 = -3.5725256e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101110010110001100010000110101;
		b = 32'b01010000010000000100001001110010;
		correct = 32'b00111111001000101100101101101011;
		#400 //4.928698e-11 * 12902320000.0 = 0.6359164
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011010111001011111001101101011;
		b = 32'b11011101010000111011110000101000;
		correct = 32'b00111000101011111101000101101101;
		#400 //-9.510544e-23 * -8.81512e+17 = 8.383659e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101011110001101010000001110100;
		b = 32'b00110010011110100110111000000111;
		correct = 32'b00011110110000100100111000010000;
		#400 //1.4113281e-12 * 1.45769325e-08 = 2.0572835e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011110100001111011110110100101;
		b = 32'b00111011101001110100011010111001;
		correct = 32'b01011010101100010110010001101101;
		#400 //4.8905777e+18 * 0.0051048663 = 2.4965745e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110001100010010101111011111101;
		b = 32'b10010001001110010010110011010100;
		correct = 32'b11000011010001101011101101100110;
		#400 //1.360457e+30 * -1.460774e-28 = -198.73203
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010101110100010111110100011011;
		b = 32'b11010010011010000010110110000100;
		correct = 32'b11101000101111011111111010011111;
		#400 //28791907000000.0 * -249299010000.0 = -7.1777936e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101111001110110100110101000011;
		b = 32'b10000000110011001100100010011110;
		correct = 32'b00110000100101011101010001011001;
		#400 //-5.79671e+28 * -1.8806409e-38 = 1.090153e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110111000111110110111101110110;
		b = 32'b01101000000000011001100000110111;
		correct = 32'b01011111101000010110101111101110;
		#400 //9.50309e-06 * 2.4479726e+24 = 2.3263304e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011010001001111000111111100010;
		b = 32'b01100000110001111101001000000110;
		correct = 32'b11111011100000101100101001010001;
		#400 //-1.179113e+16 * 1.1518862e+20 = -1.3582041e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111001101111000010001100100110;
		b = 32'b00001101110111111111000010101011;
		correct = 32'b11001000001001001001001101111101;
		#400 //-1.2210809e+35 * 1.3801375e-30 = -168525.95
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000101100001000101000011011100;
		b = 32'b11111001011101110111100001000111;
		correct = 32'b11111111011111111101000001011110;
		#400 //4234.1074 * -8.030855e+34 = -3.4003504e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001100010010000100101111010101;
		b = 32'b10111111011001101101000011011010;
		correct = 32'b11001100001101001001011110001010;
		#400 //52506452.0 * -0.9016243 = -47341096.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001111100101111111001000001011;
		b = 32'b01010001001001011101101001011100;
		correct = 32'b11100001010001001110000100111000;
		#400 //-5098444300.0 * 44520817000.0 = -2.2698691e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110101011101100001111010001000;
		b = 32'b00000011000011100111010100101101;
		correct = 32'b10111001000010001111010110010111;
		#400 //-3.1199323e+32 * 4.186456e-37 = -0.0001306146
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001010100111000011100011100001;
		b = 32'b01011100101110100000101011111101;
		correct = 32'b00100111111000110001000000010000;
		#400 //1.5043649e-32 * 4.1893142e+17 = 6.302257e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101010101100011011100010110011;
		b = 32'b11000101011010000011111100010010;
		correct = 32'b00110000101000010011101100101011;
		#400 //-3.1569677e-13 * -3715.942 = 1.1731108e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000111010100011000101101100001;
		b = 32'b01010101001001001101000000100011;
		correct = 32'b10011101000001101110011110101000;
		#400 //-1.5764372e-34 * 11325865000000.0 = -1.7854516e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110010110010000011010011000101;
		b = 32'b01000001010010111110101011001011;
		correct = 32'b11110100100111110111100101110111;
		#400 //-7.930982e+30 * 12.7448225 = -1.01078955e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010001100111011111110110110010;
		b = 32'b00011000001110000010100010111000;
		correct = 32'b00101010011000110100111011110010;
		#400 //84820770000.0 * 2.3802e-24 = 2.018904e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100000010001110100100000000100;
		b = 32'b11101001110011011000000000011111;
		correct = 32'b01001010100111111111100001100111;
		#400 //-1.6879784e-19 * -3.1054353e+25 = 5241907.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011001100000001011101011011001;
		b = 32'b10110000001001100001010110001110;
		correct = 32'b11001010001001110000011111111111;
		#400 //4529280000000000.0 * -6.042108e-10 = -2736639.8
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010010100000100011110011001001;
		b = 32'b10010010101100000111011010101111;
		correct = 32'b10100101101100111000110001010110;
		#400 //279682780000.0 * -1.1136419e-27 = -3.1146646e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111110000001101110011000010111;
		b = 32'b00011111101110111011011001011111;
		correct = 32'b11011110010001011101010001011001;
		#400 //-4.482781e+37 * 7.949929e-20 = -3.5637791e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111101101001100101000000001100;
		b = 32'b00010011000110001001011100010011;
		correct = 32'b11010001010001100100001101011001;
		#400 //-2.7633434e+37 * 1.9259583e-27 = -53220840000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011101000100101111111100011101;
		b = 32'b01000101010110011101000001001100;
		correct = 32'b10100010111110100010001110110101;
		#400 //-1.945483e-21 * 3485.0186 = -6.7800442e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000011100111000010111011100100;
		b = 32'b01111000110110101010010000000010;
		correct = 32'b01111101000001010110001111111101;
		#400 //312.36633 * 3.5476475e+34 = 1.1081656e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000011110101111110010000000101;
		b = 32'b01011111101110010011101011011110;
		correct = 32'b00100100000111000011010101101100;
		#400 //1.2688915e-36 * 2.669445e+19 = 3.3872358e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101011101010000100011101001000;
		b = 32'b11011110101001111111101100000111;
		correct = 32'b01001010110111001101011100000101;
		#400 //-1.1956902e-12 * -6.052138e+18 = 7236482.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000010010001110011101101100011;
		b = 32'b01101010101000001100110010010001;
		correct = 32'b01101101011110100100100010100100;
		#400 //49.807995 * 9.719708e+25 = 4.8411918e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000101111110000001011010101000;
		b = 32'b00111111011001110001111001100110;
		correct = 32'b00000101110111111111100111100111;
		#400 //2.333013e-35 * 0.9028076 = 2.1062619e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101010010110000101010101011110;
		b = 32'b11000100001000011000011110100101;
		correct = 32'b11101111000010001000000001010001;
		#400 //6.538278e+25 * -646.11945 = -4.2245086e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011110010110101110101010111010;
		b = 32'b10011111011001010000110001101111;
		correct = 32'b10111110010000111101111010011010;
		#400 //3.9436563e+18 * -4.850292e-20 = -0.19127885
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001101010000110101100001011000;
		b = 32'b00010001001100110110110001000110;
		correct = 32'b10011111000010001110100101100100;
		#400 //-204834180.0 * 1.4153975e-28 = -2.8992176e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101010111001001011011010010101;
		b = 32'b01010000110010000111111000100011;
		correct = 32'b00111100001100110001111101010110;
		#400 //4.0627628e-13 * 26909678000.0 = 0.010932764
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001010010001101100000001101011;
		b = 32'b01000111001101111001110001110001;
		correct = 32'b10010010000011101000110100000001;
		#400 //-9.569543e-33 * 47004.44 = -4.49811e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101011011001001010011110011000;
		b = 32'b01111010100111111101010111100010;
		correct = 32'b11100110100011101100001100100001;
		#400 //-8.1234455e-13 * 4.1495663e+35 = -3.3708777e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101011110001110110001101110100;
		b = 32'b10010100101011110100100110010001;
		correct = 32'b00000001000010001000011001001001;
		#400 //-1.4167404e-12 * -1.7699501e-26 = 2.50756e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110001000001110100100001101;
		b = 32'b11010001001100100100010001100110;
		correct = 32'b11001111111000000001101000010010;
		#400 //0.15713902 * -47853232000.0 = -7519610000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111111111101111011011000000100;
		b = 32'b10100000000001001011111100101011;
		correct = 32'b10100000100000000111001011010100;
		#400 //1.9352422 * -1.1244087e-19 = -2.176003e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000001010010100001100001101001;
		b = 32'b01100111111101110101100101011100;
		correct = 32'b11101001110000110100010000011000;
		#400 //-12.6309595 * 2.3361458e+24 = -2.9507762e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101100111011111010010110110000;
		b = 32'b01110011111010011111111101101001;
		correct = 32'b11100001010110110000110011100110;
		#400 //-6.8111836e-12 * 3.7078415e+31 = -2.525479e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100001100101110001111110110101;
		b = 32'b11100101111001010000010000100101;
		correct = 32'b11001000000001110011000111001111;
		#400 //1.0240551e-18 * -1.351873e+23 = -138439.23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010011110010011000110000101010;
		b = 32'b11010100111100000100001010000100;
		correct = 32'b10101001001111010010011111000101;
		#400 //5.0877746e-27 * -8255265000000.0 = -4.2000925e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111000011001001001011101101111;
		b = 32'b10111101110110101101011011101010;
		correct = 32'b00110110110000110110100011011100;
		#400 //-5.450047e-05 * -0.10685523 = 5.82366e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111001011011001100110101000100;
		b = 32'b01111001010010111011000011100010;
		correct = 32'b01110011001111000110101001100011;
		#400 //0.00022583181 * 6.610149e+34 = 1.492782e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000101000100001100100011110100;
		b = 32'b01110001101000100100000010011110;
		correct = 32'b11110111001101111000011101101100;
		#400 //-2316.5596 * 1.60687e+30 = -3.7224102e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111000010001101011100110111110;
		b = 32'b00111101010001000010011011000001;
		correct = 32'b01110110000110000100010001001011;
		#400 //1.6122532e+34 * 0.04788852 = 7.7208425e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100000010011001101101000000110;
		b = 32'b01101000010001101101110110010110;
		correct = 32'b01001001000111110010000111110001;
		#400 //1.735161e-19 * 3.7564644e+24 = 651807.06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110110100010010001000111010110;
		b = 32'b11100110001000110000001000101111;
		correct = 32'b11011101001011101000111100001101;
		#400 //4.0849945e-06 * -1.924465e+23 = -7.861429e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111011101010010001111010001011;
		b = 32'b01111010001000000111110110101011;
		correct = 32'b11110110010101000000110000111000;
		#400 //-0.0051611117 * 2.0832909e+35 = -1.0752097e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010101100100100000100111000111;
		b = 32'b00110100101111011000010100000000;
		correct = 32'b00001010110110000011101000101110;
		#400 //5.8984356e-26 * 3.5300764e-07 = 2.0821928e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100000101100111001111001110000;
		b = 32'b00010101010110010111010010101011;
		correct = 32'b00110110100110001001001100101001;
		#400 //1.0354324e+20 * 4.3914836e-26 = 4.5470847e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100001110000000100000101101101;
		b = 32'b00100110100010001111110001101001;
		correct = 32'b10001000110011011100000010100010;
		#400 //-1.3027744e-18 * 9.505312e-16 = -1.23832765e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000101000000111100101110010011;
		b = 32'b11100001001010000010010100110100;
		correct = 32'b10100110101011010010000101111111;
		#400 //6.196981e-36 * -1.9385836e+20 = -1.2013366e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010011110101100010110001101010;
		b = 32'b00010111010000101001100100111101;
		correct = 32'b00101011101000101100110111011100;
		#400 //1839736300000.0 * 6.2878195e-25 = 1.156793e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001100010010100011010000010111;
		b = 32'b11000000010111110110101101100000;
		correct = 32'b11001101001100000111100000110000;
		#400 //53006428.0 * -3.4909286 = -185041660.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110101110001100010111001001000;
		b = 32'b11110011111010100001100001100001;
		correct = 32'b01101010001101010011100100101101;
		#400 //-1.4765619e-06 * -3.709387e+31 = 5.4771395e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111000110010111001111010101110;
		b = 32'b10110100001101111000110011011010;
		correct = 32'b01101101100100011111111001110111;
		#400 //-3.3039208e+34 * -1.7094445e-07 = 5.6478694e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010000001100010011011000100110;
		b = 32'b01101101001000000111011111000011;
		correct = 32'b10111101110111100010100101111110;
		#400 //-3.494881e-29 * 3.103899e+27 = -0.10847758
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101001101011001111001001010111;
		b = 32'b00001100010100111100001000110101;
		correct = 32'b00110110100011110000111011110001;
		#400 //2.6134957e+25 * 1.6313291e-31 = 4.2634715e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000101111011000111000011010111;
		b = 32'b10001100111010001010111010100001;
		correct = 32'b10010011010101101110011110001100;
		#400 //7566.105 * -3.585036e-31 = -2.7124759e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011011001010000011010110110101;
		b = 32'b11001010011001101110000110110001;
		correct = 32'b10100110000101111011010010001100;
		#400 //1.3913988e-22 * -3782764.2 = -5.2633336e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010011000011110000110110100010;
		b = 32'b00101001010010100101111101111000;
		correct = 32'b00111100111000100010110000110110;
		#400 //614409040000.0 * 4.4935816e-14 = 0.027608972
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010111100000001111010101100101;
		b = 32'b10011011111000000010101111011110;
		correct = 32'b00110011111000011101100110100011;
		#400 //-283582900000000.0 * -3.708604e-22 = 1.0516967e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101000011011101111001101100100;
		b = 32'b00000001010111000101010011010100;
		correct = 32'b10101010010011011010100001011000;
		#400 //-4.513652e+24 * 4.046848e-38 = -1.8266064e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011110001000000100010101111101;
		b = 32'b01000001000111100000000110000001;
		correct = 32'b00011111110001011101011110101000;
		#400 //8.484699e-21 * 9.875367 = 8.378952e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001001111100000101101110111010;
		b = 32'b00100001010100011100001010111100;
		correct = 32'b10101011110001001111000110111001;
		#400 //-1969015.2 * 7.1069683e-19 = -1.3993729e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000100110000000110100110011;
		b = 32'b11110100000011000110011011111110;
		correct = 32'b01100101001001101100100011001000;
		#400 //-1.1063207e-09 * -4.449527e+31 = 4.9226037e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010001010000110011011111100101;
		b = 32'b01110111110110001010000001100011;
		correct = 32'b01001001101001010011000101111000;
		#400 //1.5400011e-28 * 8.787415e+33 = 1353263.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111011100011110001110011111010;
		b = 32'b01011000110111101000001101111101;
		correct = 32'b01010100111110001100100101000101;
		#400 //0.004367468 * 1957250600000000.0 = 8548229000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111011111011111010110100010010;
		b = 32'b11001000001101100000100111100101;
		correct = 32'b11000100101010100110111001001110;
		#400 //0.0073143328 * -186407.58 = -1363.447
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110010110110101110101110000100;
		b = 32'b00010000011111001001000000001001;
		correct = 32'b00000011110101111111101100000010;
		#400 //2.548564e-08 * 4.9809198e-29 = 1.2694193e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010000100110000100011000011100;
		b = 32'b01101100100100010100101000100011;
		correct = 32'b11111101101011001101011110011110;
		#400 //-20437852000.0 * 1.4051548e+27 = -2.8718345e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111101100010001011101011100000;
		b = 32'b01011010101011001100000011010001;
		correct = 32'b11011000101110001000100100010101;
		#400 //-0.066762686 * 2.431285e+16 = -1623191200000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110111001010010101100101010000;
		b = 32'b10010110110000001111011010101100;
		correct = 32'b11001110011111110100110001010011;
		#400 //3.4348033e+33 * -3.1174945e-25 = -1070798000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001110111101100010101000010011;
		b = 32'b10001001101001111001010001111010;
		correct = 32'b00011001001000010010010000111000;
		#400 //-2064976300.0 * -4.0343414e-33 = 8.330819e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100110101010001100100001000101;
		b = 32'b11111011001100010101110111100010;
		correct = 32'b01100010011010011110000010111011;
		#400 //-1.1711625e-15 * -9.209407e+35 = 1.0785712e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000001010010111010101011001000;
		b = 32'b10110111010001001001110111000010;
		correct = 32'b00111001000111000110110001000011;
		#400 //-12.729195 * -1.1719241e-05 = 0.0001491765
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100110011000001010101001010101;
		b = 32'b00100100010101001110010100001110;
		correct = 32'b00001011001110101101011000010011;
		#400 //7.7946455e-16 * 4.616419e-17 = 3.5983349e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011101101101010101111001111101;
		b = 32'b01001111100111010101001011101110;
		correct = 32'b00101101110111101110101101100111;
		#400 //4.8008e-21 * 5278915600.0 = 2.5343018e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100110100110110101000111111010;
		b = 32'b11010101000111000100100111000000;
		correct = 32'b10111100001111011010010101100110;
		#400 //1.0777505e-15 * -10740035000000.0 = -0.011575079
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101110110010101111101110000101;
		b = 32'b11110011000101001000000000010001;
		correct = 32'b01100010011010110111110111101000;
		#400 //-9.230575e-11 * -1.1765403e+31 = 1.08601434e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011100001001110000000111000100;
		b = 32'b01000100010100000001111101011001;
		correct = 32'b10100001000001111100010111100011;
		#400 //-5.5257947e-22 * 832.4898 = -4.600168e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101101100101011111011100111101;
		b = 32'b00000100001011111111011011100101;
		correct = 32'b00110010010011100010100101001001;
		#400 //5.80152e+27 * 2.068452e-36 = 1.2000165e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101010101011000101010110100000;
		b = 32'b01000001001101000100000010010101;
		correct = 32'b01101100011100101010111101011100;
		#400 //1.041698e+26 * 11.265767 = 1.17355264e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110001100101001010111000100001;
		b = 32'b10111100000100001100111010111111;
		correct = 32'b01101110001010000011010000001011;
		#400 //-1.4724573e+30 * -0.008838355 = 1.30141e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101101110011101100100010011011;
		b = 32'b11101010100111111101111000001010;
		correct = 32'b11011001000000010010000111110010;
		#400 //2.3508575e-11 * -9.663388e+25 = -2271724700000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101110100100011101011010101011;
		b = 32'b00110110000001010000110010001100;
		correct = 32'b11100101000101111001011101011001;
		#400 //-2.2567422e+28 * 1.9825848e-06 = -4.4741826e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000101111100111100111001001101;
		b = 32'b01110100110111011111001111101001;
		correct = 32'b01111011010100110110000101100011;
		#400 //7801.7876 * 1.4067928e+32 = 1.0975499e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110011011000000011110000011111;
		b = 32'b10010110101111001111111001110110;
		correct = 32'b01001010101001011000101100001010;
		#400 //-1.7765715e+31 * -3.0533626e-25 = 5424517.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000001101101001100101101110000;
		b = 32'b11100010111000111000111101101100;
		correct = 32'b01100101001000001011010110101110;
		#400 //-22.599335 * -2.0988728e+21 = 4.7433127e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110000100000101001111111010111;
		b = 32'b10011110011011010001010000111010;
		correct = 32'b01001111011100011111000010011000;
		#400 //-3.234103e+29 * -1.2550858e-20 = 4059076600.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001111110110010001001110011110;
		b = 32'b00111000011000000110100111000010;
		correct = 32'b01001000101111100100101011011000;
		#400 //7283883000.0 * 5.3504256e-05 = 389718.75
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011001100011100101010000100000;
		b = 32'b11001001000010111110101111100111;
		correct = 32'b01100011000110111001010110101010;
		#400 //-5007743000000000.0 * -573118.44 = 2.8700298e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000000111101011001011110011000;
		b = 32'b11110110010110110111101001110111;
		correct = 32'b11110111110100101000111000101011;
		#400 //7.674755 * -1.1128876e+33 = -8.5411394e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110010100101011101101101011011;
		b = 32'b10110100101001001110010000101001;
		correct = 32'b11100111110000010000110000101011;
		#400 //5.936442e+30 * -3.071339e-07 = -1.8232824e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000100101001111101011110110000;
		b = 32'b10010100011010101001011000100001;
		correct = 32'b00011001100110011100110110010101;
		#400 //-1342.7402 * -1.1843589e-26 = 1.5902863e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100111111001001111011000011011;
		b = 32'b00110111100010000001110010111100;
		correct = 32'b11011111111100110111100011100011;
		#400 //-2.1624788e+24 * 1.6225844e-05 = -3.5088044e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001110101101100110000010110010;
		b = 32'b11110100101101110011110011000000;
		correct = 32'b01000100000000101000101001100111;
		#400 //-4.495958e-30 * -1.1614044e+32 = 522.16254
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011000100101011011111110000110;
		b = 32'b01001000101111000011111101111000;
		correct = 32'b00100001110111000011101110001101;
		#400 //3.8708987e-24 * 385531.75 = 1.4923543e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010101101010000111110100100100;
		b = 32'b01001101101000101101101010111010;
		correct = 32'b01100011110101100101111001001100;
		#400 //23156929000000.0 * 341530430.0 = 7.908796e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001101011110001101110010001000;
		b = 32'b10110011001000100111101110011001;
		correct = 32'b11000001000111011111001110110101;
		#400 //260950140.0 * -3.7830976e-08 = -9.871999
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100000100001000101011011110101;
		b = 32'b01011101001000101010011100100111;
		correct = 32'b01111110001010000010101011100000;
		#400 //7.628863e+19 * 7.325237e+17 = 5.588323e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001100001110011001001111000000;
		b = 32'b00110101101000110100010110010100;
		correct = 32'b11000010011011001011011100000111;
		#400 //-48647936.0 * 1.2164696e-06 = -59.178738
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001100011100100000100101010110;
		b = 32'b11011000000011000011101100100001;
		correct = 32'b00100101000001001001010100000010;
		#400 //-1.8645811e-31 * -616742340000000.0 = 1.1499661e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110101000101001100011111111101;
		b = 32'b11110001100001011000101001010110;
		correct = 32'b11100111000110110011100010011000;
		#400 //5.542532e-07 * -1.3225198e+30 = -7.330108e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110010100110101110111101010;
		b = 32'b10101110110010100010111110100100;
		correct = 32'b10101101101001101110111101110000;
		#400 //0.20641294 * -9.194359e-11 = -1.8978347e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110000001011101100110101010000;
		b = 32'b01001011001011011101100000010010;
		correct = 32'b11111011111011010110100010010001;
		#400 //-2.163944e+29 * 11393042.0 = -2.4653904e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111110010111011110100010100001;
		b = 32'b01011111110101110110010011001101;
		correct = 32'b11011110101110101011010111000000;
		#400 //-0.21670772 * 3.1041511e+19 = -6.7269353e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110010011110111110111010001001;
		b = 32'b01011111011000110101000001000010;
		correct = 32'b01010010010111111011001101111111;
		#400 //1.46643595e-08 * 1.6379664e+19 = 240197290000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100110010101110111011010010101;
		b = 32'b00111110001110110001010010000110;
		correct = 32'b11100101000111010111010011100101;
		#400 //-2.5437406e+23 * 0.18269548 = -4.647299e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110101110100100010001011101101;
		b = 32'b10100010110000011110011001000001;
		correct = 32'b01011001000111110010100101010101;
		#400 //-5.3275914e+32 * -5.2556546e-18 = 2799998000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100011010011000010100110110000;
		b = 32'b01010010011111111110110000010100;
		correct = 32'b00110110010011000001100111001101;
		#400 //1.106769e-17 * 274794350000.0 = 3.0413387e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111100000110100010001111011000;
		b = 32'b10101001001101100010101100000111;
		correct = 32'b00100101110110110101111011001000;
		#400 //-0.00940796 * -4.044944e-14 = 3.805467e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101001100011010100111110010101;
		b = 32'b00011101010010001011001001110110;
		correct = 32'b11000111010111011001000101011110;
		#400 //-2.1354295e+25 * 2.6562042e-21 = -56721.367
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110110001101101011010111111001;
		b = 32'b00000111101110110110111111111101;
		correct = 32'b00111110100001011100011011011010;
		#400 //9.26454e+32 * 2.8202454e-34 = 0.26128274
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100111010111001110000111111001;
		b = 32'b10011000111110001110010001000010;
		correct = 32'b11000000110101101011111111011011;
		#400 //1.0430891e+24 * -6.433698e-24 = -6.71092
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001110101011111000000001110001;
		b = 32'b11010011101001000001010001111110;
		correct = 32'b01100010111000001111100010101010;
		#400 //-1472215200.0 * -1409436900000.0 = 2.0749944e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011001111111101101010000111010;
		b = 32'b11111001101011011010010010101010;
		correct = 32'b01010100001011001101100101010100;
		#400 //-2.6348702e-23 * -1.1270089e+35 = 2969522100000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011001000101011111111010111111;
		b = 32'b00001100100111010011000101101001;
		correct = 32'b00100110001110000011010001011101;
		#400 //2638741700000000.0 * 2.4219418e-31 = 6.390879e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010011011001010000001101010000;
		b = 32'b11100110101010100101111001010011;
		correct = 32'b11111010100110000110100010010101;
		#400 //983603100000.0 * -4.0227114e+23 = -3.9567515e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000001010011110100111011001011;
		b = 32'b10100010101000001010100101011101;
		correct = 32'b10100100100000100001101001100101;
		#400 //12.956737 * -4.3547407e-18 = -5.642323e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001011010110011100101010100101;
		b = 32'b11111111110010000110011101001001;
		correct = 32'b11111111110010000110011101001001;
		#400 //14273189.0 * nan = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001101010100000010111011011010;
		b = 32'b00000101011001011100010110001111;
		correct = 32'b10010011001110101101101010010001;
		#400 //-218295710.0 * 1.0803814e-35 = -2.3584262e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001101001101101111001101010100;
		b = 32'b01100000101110011000000110100110;
		correct = 32'b01101110100001001001001001111111;
		#400 //191837500.0 * 1.0693718e+20 = 2.0514562e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000011110101000011110001111110;
		b = 32'b01110001010100101110100101011011;
		correct = 32'b10110101101011101101101100010110;
		#400 //-1.2474128e-36 * 1.0443834e+30 = -1.3027773e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011001101000110001000100101000;
		b = 32'b01110010011111000011100101000010;
		correct = 32'b01001100101000001010100101011100;
		#400 //1.6860734e-23 * 4.9958043e+30 = 84232930.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000000100100100011101001111100;
		b = 32'b00011011100101111001011011000101;
		correct = 32'b00011100101011010010110100111100;
		#400 //4.569639 * 2.5078287e-22 = 1.1459872e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111101110010010001001111111101;
		b = 32'b00110100011110011110100010011111;
		correct = 32'b11110010110001000100101100101000;
		#400 //-3.3409827e+37 * 2.3274559e-07 = -7.77599e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001110011011001001010001100000;
		b = 32'b01111110110111101100100101100111;
		correct = 32'b01001101110011011110001011001011;
		#400 //2.9160686e-30 * 1.4806718e+38 = 431774050.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000001001000110101101011010100;
		b = 32'b00010010110000011001001100100010;
		correct = 32'b10010100011101110000101010111001;
		#400 //-10.209675 * 1.2216283e-27 = -1.2472428e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010100111101110111011011011011;
		b = 32'b00111110000010101010100110011111;
		correct = 32'b00010011100001100000101000001001;
		#400 //2.4987507e-26 * 0.13541268 = 3.383625e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100100010011101101010111011000;
		b = 32'b10010011110001100100000010110110;
		correct = 32'b00111000101000000010110110101110;
		#400 //-1.5261753e+22 * -5.0046037e-27 = 7.637903e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101000011110101100001111001010;
		b = 32'b10011111101001001010001001111101;
		correct = 32'b11001000101000010100010010011000;
		#400 //4.7368132e+24 * -6.9725516e-20 = -330276.75
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101011111110000010110101110101;
		b = 32'b11010110101011010100011010001000;
		correct = 32'b11000011001001111111101100011000;
		#400 //1.7634077e-12 * -95259220000000.0 = -167.98083
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010000001001011100000100101100;
		b = 32'b11000111001001000001001010101000;
		correct = 32'b01010111110101000111011110101001;
		#400 //-11123601000.0 * -42002.656 = 467220800000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110100011000110000001111000000;
		b = 32'b10111101000001001010011100110010;
		correct = 32'b11110001111010110100010001100110;
		#400 //7.1943814e+31 * -0.032386012 = -2.3299733e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100111110100010110011110110000;
		b = 32'b01100000000011101011010010111000;
		correct = 32'b01001000011010010111011010101110;
		#400 //5.812157e-15 * 4.1132185e+19 = 239066.72
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110110100011111000111110001111;
		b = 32'b00010111110101001101111100011000;
		correct = 32'b00001110111011101011111111111100;
		#400 //4.2784445e-06 * 1.3756496e-24 = 5.8856404e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101110001110010001000101111011;
		b = 32'b01100010101000111011101000111011;
		correct = 32'b01010001011011001011100110000101;
		#400 //4.2079656e-11 * 1.5101193e+21 = 63545300000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010111001001110010100111010010;
		b = 32'b01011111000011001010011001010110;
		correct = 32'b01110110101101111010111011111000;
		#400 //183798060000000.0 * 1.0134883e+19 = 1.8627717e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011011111111010010111111100111;
		b = 32'b00111100111100001000011001100001;
		correct = 32'b00011001011011011110000111010000;
		#400 //4.1886295e-22 * 0.029360952 = 1.2298215e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100100011101011011000010011001;
		b = 32'b11001001011000011010101001100111;
		correct = 32'b00101110010110001001001111000001;
		#400 //-5.327549e-17 * -924326.44 = 4.9243946e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101111011001110110100010000010;
		b = 32'b00011111111110011111101001100111;
		correct = 32'b11001111111000011111011100000000;
		#400 //-7.161738e+28 * 1.0586986e-19 = -7582122000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001001111000011010001001011011;
		b = 32'b00101111111011101010111001000101;
		correct = 32'b00111010010100100101111010001010;
		#400 //1848395.4 * 4.3415774e-10 = 0.00080249517
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000011010001000100001101001111;
		b = 32'b10100001011001010010011011101011;
		correct = 32'b10100101001011111010111000001100;
		#400 //196.26292 * -7.7639725e-19 = -1.52378e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101101001010101001100111011101;
		b = 32'b10111101100011011110000100011000;
		correct = 32'b01101011001111010001100110000000;
		#400 //-3.2999038e+27 * -0.06927699 = 2.286074e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110001011011010011011011011;
		b = 32'b11010110110100100100110011011100;
		correct = 32'b11010101100011101010011100000010;
		#400 //0.16958182 * -115613775000000.0 = -19605993000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010110101000011110100010001111;
		b = 32'b11001011000110011101001000001010;
		correct = 32'b11100010010000101001000110101001;
		#400 //89010100000000.0 * -10080778.0 = -8.972911e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101010000111001110101111011011;
		b = 32'b01001010010010111001111101100101;
		correct = 32'b00110100111110011010000101110110;
		#400 //1.3937412e-13 * 3336153.2 = 4.6497343e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000001000001101110000010111001;
		b = 32'b11111101001101100111111111001111;
		correct = 32'b01111110110000000100111000110100;
		#400 //-8.429864 * -1.5161445e+37 = 1.2780891e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010010100100111110100000111011;
		b = 32'b01100001001111111111101111110110;
		correct = 32'b11110100010111011101011110101110;
		#400 //-317628200000.0 * 2.2134274e+20 = -7.0304694e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010000000110011101011111000011;
		b = 32'b11100111001010001011111000011011;
		correct = 32'b11110111110010101100111110101101;
		#400 //10324217000.0 * -7.968644e+23 = -8.227001e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011001111011010111101000111000;
		b = 32'b10000110001001101101011011101100;
		correct = 32'b00100000100110101100010010011111;
		#400 //-8355494000000000.0 * -3.137903e-35 = 2.6218728e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110101011001100010000100101000;
		b = 32'b10110111001011101011101101100110;
		correct = 32'b11101101000111010001001011111111;
		#400 //2.9172382e+32 * -1.041484e-05 = -3.038257e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101100000110101111100111111000;
		b = 32'b10110111000110110011010001011100;
		correct = 32'b11100011101110111110101000010111;
		#400 //7.494201e+26 * -9.250911e-06 = -6.932818e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011000000000011001101110110011;
		b = 32'b11100011011011000000110001100100;
		correct = 32'b11111011111011110000001110011110;
		#400 //570022900000000.0 * -4.3543244e+21 = -2.4820646e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010010000111111111111101010000;
		b = 32'b10111001011011001011001010011100;
		correct = 32'b11001100000100111110111011111111;
		#400 //171795810000.0 * -0.00022573251 = -38779900.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110100101001000111101010100101;
		b = 32'b01000111110010110101000100011000;
		correct = 32'b10111101000000101010000101011011;
		#400 //-3.0636616e-07 * 104098.19 = -0.03189216
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101010011001111011000010001010;
		b = 32'b01111110111000101010001000010110;
		correct = 32'b11101001110011010001110010001011;
		#400 //-2.0578171e-13 * 1.5062356e+38 = -3.0995573e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101011001100000111101011110000;
		b = 32'b11010010001001001001001001001010;
		correct = 32'b01111101111000101110011100110110;
		#400 //-2.133515e+26 * -176707240000.0 = 3.7700755e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110011011111000111100101111000;
		b = 32'b10101110000100001000110010001001;
		correct = 32'b10100010000011101000111011101101;
		#400 //5.8783797e-08 * -3.286663e-11 = -1.9320253e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100011010100101000000011110101;
		b = 32'b00100110001001101010000001010111;
		correct = 32'b10001010000010010000001101110111;
		#400 //-1.14114305e-17 * 5.781012e-16 = -6.596962e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101111000111011000011110010011;
		b = 32'b10101001111010000001110111000000;
		correct = 32'b10011001100011101101010100101100;
		#400 //1.4327232e-10 * -1.03080305e-13 = -1.4768555e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001000011000110101111001001111;
		b = 32'b01001100011100111110101000111101;
		correct = 32'b11010101010110001010001010001111;
		#400 //-232825.23 * 63940852.0 = -14887043000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101011111100110011011001001110;
		b = 32'b01000100100111100110110101110010;
		correct = 32'b10110001000101101000001101111111;
		#400 //-1.7281261e-12 * 1267.4202 = -2.190262e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001101101110100000101100110010;
		b = 32'b01100100101110010110110100111000;
		correct = 32'b00110011000001101100000101110111;
		#400 //1.146583e-30 * 2.7364142e+22 = 3.137526e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110010111011101111110011000010;
		b = 32'b01100001111100100111100101100101;
		correct = 32'b01010101011000100101110001000011;
		#400 //2.7821788e-08 * 5.5910743e+20 = 15555368000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111100011011011100011101000111;
		b = 32'b10010100011011000111110011110101;
		correct = 32'b11010001010110111010011111000110;
		#400 //4.9384647e+36 * -1.19395985e-26 = -58963290000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110011001111000000011001101010;
		b = 32'b00010110111011100011110110110011;
		correct = 32'b01001010101011101111101101001000;
		#400 //1.489688e+31 * 3.8489911e-25 = 5733796.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001000111110111010000001111001;
		b = 32'b01010100010000010001010100111100;
		correct = 32'b00011101101111011100100011011010;
		#400 //1.514424e-33 * 3317139800000.0 = 5.023556e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100101010101010111010100011101;
		b = 32'b10101010110000000101000000110110;
		correct = 32'b10010000101000000101101010110111;
		#400 //1.8514485e-16 * -3.416171e-13 = -6.324864e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000111001011000001011110111110;
		b = 32'b11110011000101010101011111100001;
		correct = 32'b00111010110010001100100111001010;
		#400 //-1.2946819e-34 * -1.1832193e+31 = 0.0015318927
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100001100011000011111001101001;
		b = 32'b11100110011011101010010010101101;
		correct = 32'b11001000100000101011110000111100;
		#400 //9.503289e-19 * -2.8174024e+23 = -267745.88
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001000001010101001000101111100;
		b = 32'b01010100101010100000110100110111;
		correct = 32'b01011101011000101001101011010101;
		#400 //174661.94 * 5842929000000.0 = 1.02053735e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010000000110001101001010110001;
		b = 32'b10011010100100000110101011010101;
		correct = 32'b10101011001011000110110010010100;
		#400 //10255779000.0 * -5.97296e-23 = -6.125736e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001000011110110011001101001101;
		b = 32'b01010000111010100110101110011100;
		correct = 32'b00011001111001100000011001111100;
		#400 //7.559287e-34 * 31463367000.0 = 2.3784062e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101000011111111000011000010110;
		b = 32'b01111011101010010100111110100000;
		correct = 32'b11100100101010001111111011111111;
		#400 //-1.4184419e-14 * 1.7582263e+36 = -2.493942e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010001110000011010100111001001;
		b = 32'b00111011001010110101110001011001;
		correct = 32'b10001101100000011010001001000110;
		#400 //-3.055467e-28 * 0.0026147573 = -7.989305e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001111111001011000100110000111;
		b = 32'b11001010010001101001010110011010;
		correct = 32'b01011010101100100000111010000010;
		#400 //-7701991000.0 * -3253606.5 = 2.5059249e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000111110000010100011101110101;
		b = 32'b01001101010011110010110010100110;
		correct = 32'b00010101100111000110101001111101;
		#400 //2.908141e-34 * 217238110.0 = 6.317591e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111000000101000111111110000;
		b = 32'b00011011001101110111011011101110;
		correct = 32'b00100010101110110010001100011001;
		#400 //33423.938 * 1.5175833e-22 = 5.0723613e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000011000111010100011011100011;
		b = 32'b00110101000111111110001001000100;
		correct = 32'b10111000110001000111010000010011;
		#400 //-157.2769 * 5.9561376e-07 = -9.367629e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101001000001010100000101011101;
		b = 32'b10001110010101111100010011000111;
		correct = 32'b00110111111000001010000010100101;
		#400 //-1.0068488e+25 * -2.659554e-30 = 2.6777687e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010000100011011000110111101111;
		b = 32'b11101000000000010100011110010100;
		correct = 32'b10111001000011101111100000110011;
		#400 //5.583338e-29 * -2.4420226e+24 = -0.00013634637
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110101110000011000110010000111;
		b = 32'b00100010111010001001100110001001;
		correct = 32'b11011001001011111101101101101111;
		#400 //-4.9070485e+32 * 6.3046288e-18 = -3093712000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001010111100010000001001000111;
		b = 32'b01111100000100101011011110010010;
		correct = 32'b11000111100010100010000000011111;
		#400 //-2.3208312e-32 * 3.0471944e+36 = -70720.24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000010001001101100101001001;
		b = 32'b01000100100010010000101000010001;
		correct = 32'b10110101010100101100000000001011;
		#400 //-7.1613165e-10 * 1096.3146 = -7.8510556e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101100100100001010111100101000;
		b = 32'b00100101011010110101101000101101;
		correct = 32'b01010010100001010000001111000001;
		#400 //1.3992998e+27 * 2.0413554e-16 = 285646800000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010000111001101010111010001100;
		b = 32'b00011110000111011001011000011010;
		correct = 32'b10101111100011100000000001001110;
		#400 //-30961590000.0 * 8.342551e-21 = -2.5829866e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010001101001001111001111101100;
		b = 32'b01010000001110101101101101100001;
		correct = 32'b00100010011100001100110100101001;
		#400 //2.6024966e-28 * 12539758000.0 = 3.2634676e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100111011011111110011000011010;
		b = 32'b11011000010100011001000101001011;
		correct = 32'b11000000010001000110001100000011;
		#400 //3.3292651e-15 * -921687840000000.0 = -3.0685432
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101000100000111111111010101010;
		b = 32'b01001000001110110101110001001010;
		correct = 32'b01110001010000010011010100111000;
		#400 //4.986622e+24 * 191857.16 = 9.567191e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111111110001101011110101110111;
		b = 32'b00011010001101001101011011110000;
		correct = 32'b00011010100011000110010000010100;
		#400 //1.552657 * 3.7396753e-23 = 5.806433e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011001001001011100000011001000;
		b = 32'b10101011010011001001010111011000;
		correct = 32'b11000101000001000111011010100100;
		#400 //2915958500000000.0 * -7.268331e-13 = -2119.415
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111101100111100111011110010101;
		b = 32'b10011011110001100100111001010011;
		correct = 32'b11011001111101011000000111110010;
		#400 //2.6329866e+37 * -3.2806968e-22 = -8638030700000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111101000011110100011100001010;
		b = 32'b00101001010110001001101100011011;
		correct = 32'b11100110111100100111010101111111;
		#400 //-1.1903029e+37 * 4.8096167e-14 = -5.7249005e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010111011110011110101110110111;
		b = 32'b00010110001010110110101111101000;
		correct = 32'b10101110001001110101100111001011;
		#400 //-274790780000000.0 * 1.3847319e-25 = -3.8051156e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011100001001011000110011011101;
		b = 32'b01001100001100111011110010110110;
		correct = 32'b11101000111010000111011100001111;
		#400 //-1.86393e+17 * 47117016.0 = -8.782282e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010011001011101011100010111000;
		b = 32'b01000001011001111100101011101000;
		correct = 32'b00010101000111100011001100101010;
		#400 //2.2052961e-27 * 14.487038 = 3.1948207e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101111001110101000011100101111;
		b = 32'b01101000010011100100100101100010;
		correct = 32'b11011000000101100100111001000000;
		#400 //-1.6964628e-10 * 3.8966447e+24 = -661051300000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111101101100111101111010010100;
		b = 32'b00001000000010101100011001111101;
		correct = 32'b10000110010000110000001011100100;
		#400 //-0.08782688 * 4.1761186e-34 = -3.6677547e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100110011110010100001100100110;
		b = 32'b10011001110000010100011011100101;
		correct = 32'b01000000101111000011000010100111;
		#400 //-2.9427698e+23 * -1.9984366e-23 = 5.880939
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100001000000100111101100111001;
		b = 32'b10100011100101001111001001000010;
		correct = 32'b11000101000101111101010101101110;
		#400 //1.5043474e+20 * -1.6148792e-17 = -2429.3394
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000011101111001000001111011111;
		b = 32'b00111110011000111001010010010000;
		correct = 32'b00000010101001111001011001010101;
		#400 //1.1079923e-36 * 0.22224641 = 2.462473e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110110010011101011110000000101;
		b = 32'b01001000000011011111001011010010;
		correct = 32'b11111110111001010100001101001100;
		#400 //-1.0482682e+33 * 145355.28 = -1.5237132e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111011101100111111100001000001;
		b = 32'b01001011110001000010111000011011;
		correct = 32'b01001000000010011110101001111011;
		#400 //0.0054922407 * 25713718.0 = 141225.92
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001000101001000000101011011101;
		b = 32'b01101101111010110110111000101010;
		correct = 32'b01110111000101101101110010010000;
		#400 //335958.9 * 9.1077697e+27 = 3.0598362e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101000010011110101001100110011;
		b = 32'b00011011001001101110001010000001;
		correct = 32'b01000100000001110010011101100011;
		#400 //3.9162585e+24 * 1.3804386e-22 = 540.6154
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000011100101010100110111000111;
		b = 32'b00001011010110111011100100101011;
		correct = 32'b00001111100000000010010110001000;
		#400 //298.60764 * 4.231717e-32 = 1.2636231e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111000011111011100110011111010;
		b = 32'b00001000110011110010111111001001;
		correct = 32'b10000001110011010110100000011110;
		#400 //-6.05108e-05 * 1.2469594e-33 = -7.545451e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100001111100101011110011111111;
		b = 32'b11100101000111110000011101010110;
		correct = 32'b01000111100101101100101001010111;
		#400 //-1.6448585e-18 * -4.6936975e+22 = 77204.68
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001001000110110000011110011100;
		b = 32'b11000110111000101011010110111000;
		correct = 32'b11010000100010010100101011000100;
		#400 //635001.75 * -29018.86 = -18427027000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111101001100010110011010010001;
		b = 32'b00101111110101011010011011111111;
		correct = 32'b11101101100101000000111000010000;
		#400 //-1.473787e+37 * 3.8863132e-10 = -5.727598e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001001000001000011011000110010;
		b = 32'b11100110000001101101101000100011;
		correct = 32'b00101111100010110100101000001101;
		#400 //-1.5914405e-33 * -1.5920526e+23 = 2.533657e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010000101100101011111010100010;
		b = 32'b10101001111000011110100001001010;
		correct = 32'b00111011000111011011101110111101;
		#400 //-23990702000.0 * -1.0032303e-13 = 0.00240682
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011000111100101001101100100011;
		b = 32'b11001010001010110100100000111101;
		correct = 32'b10100011101000100101001000010110;
		#400 //6.271218e-24 * -2806287.2 = -1.759884e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111111111100101000110101000110;
		b = 32'b11000001110110001101110110100010;
		correct = 32'b11000010010011010111100100110001;
		#400 //1.8949363 * -27.10822 = -51.36835
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011011100110001011001011100010;
		b = 32'b10100101011001010000100000010110;
		correct = 32'b10000001100010001001110011010111;
		#400 //2.526189e-22 * -1.9865323e-16 = -5.0183564e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011010100100111100111100111010;
		b = 32'b01111001010100000010110101011011;
		correct = 32'b01010100011100000110010100011110;
		#400 //6.113257e-23 * 6.7557354e+34 = 4129954500000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010011010101110011110110101011;
		b = 32'b01110010011000000011100101101001;
		correct = 32'b01000110001111001000011000111011;
		#400 //2.716722e-27 * 4.441219e+30 = 12065.558
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001000101110001111000001101111;
		b = 32'b11011111001110100110000000100011;
		correct = 32'b10101000100001101010010000100100;
		#400 //1.1130623e-33 * -1.3429773e+19 = -1.4948173e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100011001010010101100101001110;
		b = 32'b00100110000001101100000011111001;
		correct = 32'b01001001101100100100100011001101;
		#400 //3.1239348e+21 * 4.6752116e-16 = 1460505.6
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011001100101001010101001010011;
		b = 32'b10101010111001101011001100000011;
		correct = 32'b00000101000001011111100011111011;
		#400 //-1.5371635e-23 * -4.0980422e-13 = 6.2993604e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110011001011110001100001101000;
		b = 32'b10010010100000111100110010010111;
		correct = 32'b01000110001101000100101011011000;
		#400 //-1.3872482e+31 * -8.317698e-28 = 11538.711
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110011100010010111010011011100;
		b = 32'b10101101011111000110011001100001;
		correct = 32'b01100001100001111000011000000001;
		#400 //-2.178085e+31 * -1.4347274e-11 = 3.124958e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000010000101000100010111101011;
		b = 32'b11010001011010000010100110001100;
		correct = 32'b01010100000001100111011101101101;
		#400 //-37.06828 * -62320590000.0 = 2310117000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101010011011011100111111111101;
		b = 32'b10110111001101111100011000010011;
		correct = 32'b00100010001010101011011110101110;
		#400 //-2.1121989e-13 * -1.0953768e-05 = 2.3136535e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011110100100001001111110111101;
		b = 32'b11001110100101111111001111011111;
		correct = 32'b10101101101010111010111111111100;
		#400 //1.531266e-20 * -1274671000.0 = -1.9518602e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110000001110111000000100101100;
		b = 32'b01001110010011000100000101011100;
		correct = 32'b01111111000101011001101011001110;
		#400 //2.3211942e+29 * 856708860.0 = 1.9885876e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101111000100110011110010111110;
		b = 32'b01101101011110101111001110000010;
		correct = 32'b01011101000100000101010101011111;
		#400 //1.3391152e-10 * 4.8541022e+27 = 6.500202e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011101011111000000000011010100;
		b = 32'b10011001101111110111000100100101;
		correct = 32'b00110111101111000111001111111111;
		#400 //-1.1349217e+18 * -1.9794636e-23 = 2.2465361e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001010000011001110001010001011;
		b = 32'b11010011001001100100001011110000;
		correct = 32'b10011101101101101111111101111001;
		#400 //6.783363e-33 * -714087600000.0 = -4.843915e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111100100001010110000111000100;
		b = 32'b11000010001000110011000100100111;
		correct = 32'b11111111001010100000110110111000;
		#400 //5.540467e+36 * -40.798 = -2.2604e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011001111010111011111001110110;
		b = 32'b00111101011110001000000011010101;
		correct = 32'b00010111111001001101011100100110;
		#400 //2.4375357e-23 * 0.06066974 = 1.4788466e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011101101000101000011100110101;
		b = 32'b11011011100101000011100101101011;
		correct = 32'b01111001101111000011010100111101;
		#400 //-1.4639235e+18 * -8.344286e+16 = 1.2215395e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101110110010101011011010000001;
		b = 32'b00011011110000101000111111010000;
		correct = 32'b00001011000110100001000000101110;
		#400 //9.218316e-11 * 3.2187544e-22 = 2.9671493e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100001100000011010001111100011;
		b = 32'b00011111011011000100001110100010;
		correct = 32'b10000001011011110100101010101010;
		#400 //-8.78476e-19 * 5.003089e-20 = -4.3950936e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010110001001101011000001010101;
		b = 32'b01000010010100101000001100100011;
		correct = 32'b11011001000010010001001000001001;
		#400 //-45819068000000.0 * 52.628063 = -2411368900000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100010111011001101110000110111;
		b = 32'b11100110110111011110111011101000;
		correct = 32'b11001010010011010101011100100111;
		#400 //6.420109e-18 * -5.24025e+23 = -3364297.8
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000011000111100001111000101010;
		b = 32'b01001000100000010110100111001111;
		correct = 32'b10001100000111111101110100011011;
		#400 //-4.6466654e-37 * 265038.47 = -1.2315451e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111010101101100001101111101001;
		b = 32'b11110011011111001000100110000001;
		correct = 32'b11101110101100111010010101001010;
		#400 //0.0013893816 * -2.0008052e+31 = -2.779882e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110100010111010100000010100101;
		b = 32'b10010101010110100101000000011001;
		correct = 32'b00001010001111001010111001000110;
		#400 //-2.0605746e-07 * -4.4087935e-26 = 9.084648e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111010011000101101110101111100;
		b = 32'b10001111111001001111111000101101;
		correct = 32'b10001010110010101110111010000010;
		#400 //0.00086542196 * -2.258044e-29 = -1.9541609e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111011110010100000100111101110;
		b = 32'b10001011110110010011011000001011;
		correct = 32'b00001000001010110110110100010010;
		#400 //-0.0061657345 * -8.3666674e-32 = 5.158665e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011001010111011000100000111101;
		b = 32'b00001011010000101000010010100111;
		correct = 32'b10100101001010000101010000001001;
		#400 //-3897235300000000.0 * 3.7462837e-32 = -1.460015e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101010010100111110000100101111;
		b = 32'b00111000001010010101000111101100;
		correct = 32'b00100011000011000010001101110110;
		#400 //1.8818691e-13 * 4.0369036e-05 = 7.596924e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111101111100010000111101110100;
		b = 32'b01010000111010000011110111111100;
		correct = 32'b11001111010110101011000001011111;
		#400 //-0.117705256 * 31171010000.0 = -3668991700.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101101011101110010001001110000;
		b = 32'b11000111110100111010010011000111;
		correct = 32'b10110101110011000101000001110100;
		#400 //1.4047971e-11 * -108361.555 = -1.5222599e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000011001110110000001011100000;
		b = 32'b00011101100111101110100100111011;
		correct = 32'b10100001011010000010110001001110;
		#400 //-187.01123 * 4.2063406e-21 = -7.8663294e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100010000011000110110000101010;
		b = 32'b10011001111100101111000001010001;
		correct = 32'b10111100100001010100001000010010;
		#400 //6.4758455e+20 * -2.5119277e-23 = -0.016266856
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000000010111110110111111110011;
		b = 32'b00001000101110011101001111110001;
		correct = 32'b00001001101000100011000011100010;
		#400 //3.4912078 * 1.118411e-33 = 3.904605e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001011110111010010001000001010;
		b = 32'b10001100111001101000111101110100;
		correct = 32'b10011001010001110010100001111111;
		#400 //28984340.0 * -3.5523449e-31 = -1.0296237e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000001001101000011100000100000;
		b = 32'b01001101111000001000001011011111;
		correct = 32'b01001111100111100000110100111101;
		#400 //11.263702 * 470834140.0 = 5303335400.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110010010000010110110111111;
		b = 32'b11110101000100010001111010010101;
		correct = 32'b01101011111000101111001110100110;
		#400 //-2.982895e-06 * -1.8396077e+32 = 5.4873566e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000001000010101101111000001110;
		b = 32'b10011001101111010100111000111110;
		correct = 32'b10011011010011010110000011000011;
		#400 //8.679213 * -1.9573744e-23 = -1.6988468e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010011111101010100001001110011;
		b = 32'b01010110000101001000100010010011;
		correct = 32'b00101010100011100100110101000011;
		#400 //6.191222e-27 * 40828576000000.0 = 2.5277878e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000011011111001001000011111111;
		b = 32'b00111100101101110111000000000001;
		correct = 32'b10000000101101001111101000100111;
		#400 //-7.422259e-37 * 0.022392275 = -1.6620127e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111101100111011101011000110100;
		b = 32'b00010011101101101111000011000101;
		correct = 32'b11010001111000011001010101110110;
		#400 //-2.6225125e+37 * 4.6180676e-27 = -121109400000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110101111010111010100000011100;
		b = 32'b11101000111100000010100111010010;
		correct = 32'b01011111010111010001010000011001;
		#400 //-1.7557791e-06 * -9.073115e+24 = 1.5930385e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100101101111111010010111111111;
		b = 32'b01100111110100001001101001111010;
		correct = 32'b01001110000111000010101010000100;
		#400 //3.3245702e-16 * 1.9702036e+24 = 655008000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100001100011111011011101101111;
		b = 32'b10101001000001010001100011111011;
		correct = 32'b10001011000101010111000010100110;
		#400 //9.738611e-19 * -2.95536e-14 = -2.8781103e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011001010010010101000001111110;
		b = 32'b01010001000000110111101001011001;
		correct = 32'b11101010110011101100100011001110;
		#400 //-3541560800000000.0 * 35293336000.0 = -1.249935e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000011101001001111110111000101;
		b = 32'b10110011001110011000100001111001;
		correct = 32'b00110111011011110010011010110000;
		#400 //-329.98257 * -4.319779e-08 = 1.4254518e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110100100000110000111001111011;
		b = 32'b00010001011010010111001100101110;
		correct = 32'b11000110011011110000011001001010;
		#400 //-8.306697e+31 * 1.8415952e-28 = -15297.572
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010011001110011001101001010011;
		b = 32'b11011001100101110010010111101101;
		correct = 32'b10101101010110110010101100001100;
		#400 //2.342637e-27 * -5318052700000000.0 = -1.2458267e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100011111010101010100001011110;
		b = 32'b10101100101110011011010011101011;
		correct = 32'b01010001001010100011100110000010;
		#400 //-8.6573405e+21 * -5.278102e-12 = 45694330000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001001100011111001010100111110;
		b = 32'b11110010010100001111100010111100;
		correct = 32'b00111100011010100110100110001001;
		#400 //-3.4566344e-33 * -4.1391093e+30 = 0.014307388
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110110010111101111000001110100;
		b = 32'b10110100001011100001110100011110;
		correct = 32'b11101011000101111010000011001010;
		#400 //1.1304364e+33 * -1.6215606e-07 = -1.833071e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001111110001010010111101000111;
		b = 32'b01100101100010010000101110001100;
		correct = 32'b00110101110100110001111001100100;
		#400 //1.944391e-29 * 8.089715e+22 = 1.572957e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000101011111010000001101010;
		b = 32'b10010100001010110100111010110100;
		correct = 32'b00000101011010110000110001001010;
		#400 //-1.2778518e-09 * -8.648815e-27 = 1.1051904e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110100100111101111010000111010;
		b = 32'b00010001000110111011101000011100;
		correct = 32'b11000110010000010110001011011100;
		#400 //-1.0074907e+32 * 1.2284693e-28 = -12376.715
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001100001111001110001111110000;
		b = 32'b01000010101010000110011101000111;
		correct = 32'b01001111011110001000001110010011;
		#400 //49516480.0 * 84.20171 = 4169372400.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001100111000101000111100011000;
		b = 32'b01000111000001101100100111011101;
		correct = 32'b00010100011011101001001100011001;
		#400 //3.4906935e-31 * 34505.863 = 1.2044939e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100010111001000101101011011000;
		b = 32'b00110101001100110010001010001101;
		correct = 32'b11011000100111111100101001010111;
		#400 //-2.1062018e+21 * 6.6732974e-07 = -1405531100000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011100010100110001111001101011;
		b = 32'b00010110110000001100100011010001;
		correct = 32'b10110011100111101111110001101100;
		#400 //-2.3769866e+17 * 3.1146006e-25 = -7.4033636e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011011011001001010100101001010;
		b = 32'b01000111111011111111100101001100;
		correct = 32'b10100011110101100101100010111001;
		#400 //-1.8914418e-22 * 122866.59 = -2.3239502e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101111010101001000101011011101;
		b = 32'b00101001110100010111110101001101;
		correct = 32'b10011001101011011110110101100110;
		#400 //-1.9330622e-10 * 9.303201e-14 = -1.7983665e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100000010100001110010001101110;
		b = 32'b01100011100010110001101010110111;
		correct = 32'b11000100011000110000001110101001;
		#400 //-1.7693866e-19 * 5.132045e+21 = -908.0572
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000010100011011101101010100101;
		b = 32'b01111001001111100011110101000000;
		correct = 32'b00111100010100101101010001101110;
		#400 //2.0843584e-37 * 6.173617e+34 = 0.01286803
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011001110010010000110110100001;
		b = 32'b10101001110101011001110000101111;
		correct = 32'b11000100001001111100001100000000;
		#400 //7073932000000000.0 * -9.486194e-14 = -671.0469
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001110010111000010110011000111;
		b = 32'b01000001101100001011011110111101;
		correct = 32'b00010000100101111111110011001111;
		#400 //2.7138653e-30 * 22.089716 = 5.994851e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000110001010111111011010110100;
		b = 32'b10101100101000000111101010000101;
		correct = 32'b00110011010101111001100011111011;
		#400 //-11005.676 * -4.561076e-12 = 5.0197723e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010011100110110100010000010001;
		b = 32'b00101111111001001011000001101110;
		correct = 32'b01000100000010101011001110100001;
		#400 //1333723800000.0 * 4.159832e-10 = 554.8067
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000111011111100110011110100100;
		b = 32'b00110001111111001101101000111000;
		correct = 32'b10111001111110110100011011100001;
		#400 //-65127.64 * 7.358974e-09 = -0.0004792726
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111101111000011111001001001100;
		b = 32'b00000111110000110101000111110101;
		correct = 32'b00000110001011000110001111100110;
		#400 //0.110325426 * 2.938851e-34 = 3.2422998e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101111100010000010110010100000;
		b = 32'b10011110111101111110100100001100;
		correct = 32'b01001111000000111101111100000101;
		#400 //-8.428782e+28 * -2.6248528e-20 = 2212431000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100101000101010101010011011100;
		b = 32'b11110000010110000100100010011100;
		correct = 32'b01010101111111000101001111101001;
		#400 //-1.2952441e-16 * -2.6774617e+29 = 34679665000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000110001110000011101110110101;
		b = 32'b11000100001001011100000100110000;
		correct = 32'b01001010111011101001001100000110;
		#400 //-11790.927 * -663.01855 = 7817603.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110000010100010001001111001;
		b = 32'b01111000011100011000001001100100;
		correct = 32'b01110111000000100101000011001111;
		#400 //0.13489713 * 1.9593565e+34 = 2.6431156e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110001000010010100100101010111;
		b = 32'b10010101011001111001001011010010;
		correct = 32'b11000110111110000101111111010100;
		#400 //6.7980974e+29 * -4.67659e-26 = -31791.914
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111100011011111100101000111110;
		b = 32'b11101011001010010100101001110110;
		correct = 32'b11101000000111101001001001000010;
		#400 //0.014635621 * -2.046601e+26 = -2.9953275e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101111101100000011101111111110;
		b = 32'b01000001110011011011000100010011;
		correct = 32'b00110010000011011001100111110001;
		#400 //3.205684e-10 * 25.711462 = 8.242282e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000110111011001001110011111001;
		b = 32'b00010110011101001001100110110010;
		correct = 32'b00011101111000100001001110101100;
		#400 //30286.486 * 1.9758661e-25 = 5.9842042e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101001110100001110100100100100;
		b = 32'b00100100011010110000101000111111;
		correct = 32'b01001110101111111100111001100001;
		#400 //3.1569693e+25 * 5.096618e-17 = 1608986800.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100010101111101110110001001010;
		b = 32'b00000111110001000000011001000110;
		correct = 32'b10101011000100100011000110010110;
		#400 //-1.7609539e+21 * 2.949449e-34 = -5.1938434e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001000011101111010001100110000;
		b = 32'b01010001100111111000000000111110;
		correct = 32'b01011010100110100100101001101000;
		#400 //253580.75 * 85631420000.0 = 2.1714478e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101011001111000001100001011010;
		b = 32'b00001100011100111101000101010001;
		correct = 32'b00111000001100110010010011101001;
		#400 //2.2739305e+26 * 1.8783028e-31 = 4.27113e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101101100010001001000111111110;
		b = 32'b10101000101000000010101101010011;
		correct = 32'b00010110101010101110010010110111;
		#400 //-1.5526243e-11 * -1.7782357e-14 = 2.760932e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101010110010010010100011010100;
		b = 32'b11010111011101100100111010011101;
		correct = 32'b11000010110000011000101100000010;
		#400 //3.5733103e-13 * -270817500000000.0 = -96.7715
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111100100000001100111001101011;
		b = 32'b00100101001001110011011000001111;
		correct = 32'b00100010001010000100001110110110;
		#400 //0.015723428 * 1.4503257e-16 = 2.2804091e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111101010111110010111100101010;
		b = 32'b10011111001010010000100000101010;
		correct = 32'b10011101000100110101110101000001;
		#400 //0.05448834 * -3.5793895e-20 = -1.95035e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010110101000110111110011011010;
		b = 32'b11010100000010100101010011001111;
		correct = 32'b11101011001100001010111011101101;
		#400 //89878314000000.0 * -2376513400000.0 = -2.13597e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001100110010011001100000001000;
		b = 32'b10110110111000101010000100110111;
		correct = 32'b00000100001100100111011100101011;
		#400 //-3.1060454e-31 * -6.7540927e-06 = 2.0978519e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000101000110111000001110101001;
		b = 32'b10110100011000011111010101010000;
		correct = 32'b10111010000010010100001110111101;
		#400 //2488.2288 * -2.1044002e-07 = -0.0005236229
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101111101010000100010100101100;
		b = 32'b10011000011100101001111000111000;
		correct = 32'b10001000100111110111100101100011;
		#400 //3.0608172e-10 * -3.1357647e-24 = -9.598002e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000100011011000000011001001000;
		b = 32'b01000110111011000010101000000011;
		correct = 32'b00001011110110011011110010000110;
		#400 //2.774455e-36 * 30229.006 = 8.386902e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010110111101010011001101010010;
		b = 32'b11110010011100001111000001101001;
		correct = 32'b11001001111001101100011001100010;
		#400 //3.9614272e-25 * -4.7722906e+30 = -1890508.2
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001110111000010111000100000001;
		b = 32'b00111000111001110111100001110011;
		correct = 32'b00001000010010111101011100001010;
		#400 //5.55756e-30 * 0.00011037374 = 6.1340868e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001000001100100100100010000100;
		b = 32'b00110100010000011101100000010110;
		correct = 32'b00111101000001101111111100101000;
		#400 //182562.06 * 1.8053137e-07 = 0.03295818
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011111110101100111100110101001;
		b = 32'b10111111110101000010101001011101;
		correct = 32'b11100000001100011100000000111110;
		#400 //3.0909139e+19 * -1.6575428 = -5.123322e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010110000110011101100101000001;
		b = 32'b01010100011110100001000001011010;
		correct = 32'b01101011000101100100011111111101;
		#400 //42289594000000.0 * 4296064600000.0 = 1.8167883e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101111000001110101010000010001;
		b = 32'b01101001111001111111101101111110;
		correct = 32'b01011001011101010100001110011011;
		#400 //1.2308045e-10 * 3.5056188e+25 = 4314731400000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001011101010000111111001100101;
		b = 32'b10100101000001001001000011001111;
		correct = 32'b10110001001011101000000011110111;
		#400 //22084810.0 * -1.1498238e-16 = -2.539364e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110011110010001100111011001011;
		b = 32'b00011111110001111110010000000111;
		correct = 32'b11010100000111001100101110011101;
		#400 //-3.1819264e+31 * 8.465702e-20 = -2693723800000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001011001100101110100101000100;
		b = 32'b01011000010000001111000011011111;
		correct = 32'b01100100000001101101011101001010;
		#400 //11725124.0 * 848563060000000.0 = 9.949508e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110010110000001010101000100010;
		b = 32'b00110000110011110111010001101101;
		correct = 32'b00100100000111000010000100110001;
		#400 //2.242911e-08 * 1.5094322e-09 = 3.3855222e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000111001010101000110000001001;
		b = 32'b11111110100001111001110111001111;
		correct = 32'b11000110001101001011000111110101;
		#400 //1.2830531e-34 * -9.013258e+37 = -11564.489
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001100101110001100010011010010;
		b = 32'b10110011000011000110110000110000;
		correct = 32'b11000000010010101011001101110001;
		#400 //96872080.0 * -3.2694686e-08 = -3.1672022
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101011111101100011101100100001;
		b = 32'b00100001001000001111110011000010;
		correct = 32'b11001101100110101101100000010001;
		#400 //-5.9534996e+26 * 5.454463e-19 = -324731420.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100110000110010000001101000101;
		b = 32'b10101111101011110001011101101001;
		correct = 32'b11010110010100010100111001110100;
		#400 //1.806456e+23 * -3.1848948e-10 = -57533720000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100100100101111110100001000101;
		b = 32'b10011010111101111110110100100000;
		correct = 32'b11000000000100110001110111010000;
		#400 //2.241756e+22 * -1.025399e-22 = -2.2986946
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011110010111010011111000101010;
		b = 32'b01001111010101011000100101111011;
		correct = 32'b00101110001110001000101110001010;
		#400 //1.1712498e-20 * 3582557000.0 = 4.1960692e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011111011010010011110001011001;
		b = 32'b01001011100011010100011011110001;
		correct = 32'b01101011100000001011011011011111;
		#400 //1.6806406e+19 * 18517474.0 = 3.1121218e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101101000011111100010100101110;
		b = 32'b10001010010101111111111101011100;
		correct = 32'b10110111111100101001110000000101;
		#400 //2.7809208e+27 * -1.0399901e-32 = -2.89213e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011110010000011111110011110101;
		b = 32'b11001010011010111100111101001101;
		correct = 32'b11101001001100101011000001001011;
		#400 //3.4945792e+18 * -3863507.2 = -1.3501332e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010100111011011101000111011010;
		b = 32'b11000100001011000111011000010001;
		correct = 32'b01011001101000000011011010101101;
		#400 //-8171424000000.0 * -689.8448 = 5637014000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001010111011101001011110001111;
		b = 32'b10110000011100000001001100001001;
		correct = 32'b10111011110111111011111111010100;
		#400 //7818183.5 * -8.733854e-10 = -0.0068282876
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001000110111000000111111011000;
		b = 32'b11010100001110101111011110010111;
		correct = 32'b01011101101000001011100001011000;
		#400 //-450686.75 * -3212071100000.0 = 1.4476379e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010100011110110110111110001100;
		b = 32'b11010101000011111011100111101101;
		correct = 32'b01101010000011010010100111101100;
		#400 //-4319633000000.0 * -9876794000000.0 = 4.266413e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010001100000011101111100100010;
		b = 32'b01101001011110010011110101000111;
		correct = 32'b11111011011111001110001000111101;
		#400 //-69724290000.0 * 1.8831994e+25 = -1.3130475e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110010111100001000110101101101;
		b = 32'b00001111100101010011100011000110;
		correct = 32'b00000011000011000011011110101001;
		#400 //2.800399e-08 * 1.4714403e-29 = 4.1206197e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010101001100110001010001111101;
		b = 32'b01000101000100001000111101010010;
		correct = 32'b10011010110010100011111110010000;
		#400 //-3.6164925e-26 * 2312.9575 = -8.364793e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111000010001001110011110110001;
		b = 32'b11110011010011100001011111110100;
		correct = 32'b01101100000111101000010011011101;
		#400 //-4.694582e-05 * -1.6328415e+31 = 7.665508e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100000000101101110100100011111;
		b = 32'b00101111110000110011010011100011;
		correct = 32'b10010000011001100010010110000000;
		#400 //-1.2782628e-19 * 3.5507872e-10 = -4.538839e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100101100000100010000010110110;
		b = 32'b10010000100100110101001011010010;
		correct = 32'b00110110100101011100010111000011;
		#400 //-7.681388e+22 * -5.810888e-29 = 4.4635685e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010110100011001010101111110;
		b = 32'b00111011010100011011110000000111;
		correct = 32'b10110110101010111011010011111011;
		#400 //-0.0015989987 * 0.0032002942 = -5.117266e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111000001110000101100101101110;
		b = 32'b10101000101000110101001100110000;
		correct = 32'b01100001011010110011100110110001;
		#400 //-1.4956195e+34 * -1.8132712e-14 = 2.7119637e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001001011010010011110111001111;
		b = 32'b01111110100111101100001011011000;
		correct = 32'b11001000100100001010010110101011;
		#400 //-2.8075417e-33 * 1.0551485e+38 = -296237.34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101001010001111010010011001011;
		b = 32'b01101100100110001001001111001110;
		correct = 32'b11010110011011011111101000111010;
		#400 //-4.432981e-14 * 1.4756377e+27 = -65414743000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111011011110001100101001011100;
		b = 32'b11111000111110101100010011111011;
		correct = 32'b01110100111100111011010100001101;
		#400 //-0.0037962412 * -4.068967e+34 = 1.5446781e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111000011011111100111101111001;
		b = 32'b00001010001111011011101111100100;
		correct = 32'b11000011001100011011110000101110;
		#400 //-1.9455734e+34 * 9.135357e-33 = -177.73508
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000010010001111101110000110100;
		b = 32'b01111000110111110101111101000010;
		correct = 32'b10111011101011100110001100110000;
		#400 //-1.4683406e-37 * 3.6244196e+34 = -0.0053218827
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110001000100000110110011111110;
		b = 32'b01000011000110100010111001100100;
		correct = 32'b10110100101011011111011101111010;
		#400 //-2.1016713e-09 * 154.18121 = -3.2403824e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010100101010100111110100010010;
		b = 32'b11110110100100011011110000001000;
		correct = 32'b11001011110000100001110000100001;
		#400 //1.7214945e-26 * -1.4779234e+33 = -25442370.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001101100111100000010011010000;
		b = 32'b10101110001111011110001000010101;
		correct = 32'b10111100011010100110101000110110;
		#400 //331389440.0 * -4.3174426e-11 = -0.014307549
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110000111001011110010000110111;
		b = 32'b11000111111110001100101011000111;
		correct = 32'b10111001010111110110101100101110;
		#400 //1.6726805e-09 * -127381.555 = -0.00021306865
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111010100011101011010000110011;
		b = 32'b10110111010001001000010011100100;
		correct = 32'b01110010010110110001100000010110;
		#400 //-3.704805e+35 * -1.1713451e-05 = 4.3396055e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110001000001101111010111100;
		b = 32'b10000010110011010000111111000011;
		correct = 32'b10000001100000001101110001000100;
		#400 //0.15709966 * -3.013109e-37 = -4.733584e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011100001000110111101010000011;
		b = 32'b01100000001100010110001110011010;
		correct = 32'b11111100111000101000111010011111;
		#400 //-1.840605e+17 * 5.112892e+19 = -9.410814e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110101001001111110011001000000;
		b = 32'b00111111110000011110010111010111;
		correct = 32'b11110101011111100101011010101000;
		#400 //-2.128378e+32 * 1.5148267 = -3.2241235e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101011010101110111101110010111;
		b = 32'b00011001001010011000100001101110;
		correct = 32'b10000101000011101011001101101101;
		#400 //-7.655486e-13 * 8.764647e-24 = -6.709763e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111001111011011100110010100111;
		b = 32'b00011100100111011110001010000011;
		correct = 32'b10010111000100101010100011101011;
		#400 //-0.0004535664 * 1.044794e-21 = -4.738835e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100111011001011000101101010001;
		b = 32'b00000101011110010011101001100110;
		correct = 32'b10101101010111110111100011011111;
		#400 //-1.08399186e+24 * 1.171865e-35 = -1.2702921e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111110100000001100001010000001;
		b = 32'b00100011010111010100111101101110;
		correct = 32'b10100010010111101001111110111001;
		#400 //-0.25148395 * 1.1997254e-17 = -3.0171167e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001111100010000000010000001111;
		b = 32'b10100001001011101100001110111101;
		correct = 32'b00110001001110011011010110000011;
		#400 //-4563934700.0 * -5.921255e-19 = 2.702422e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010011010110011011101111000110;
		b = 32'b11010000001110001111111011011010;
		correct = 32'b10100100000111010101011110111000;
		#400 //2.748183e-27 * -12414839000.0 = -3.411825e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110111010100001100000100110001;
		b = 32'b00101000000110011010110001101001;
		correct = 32'b01011111111110101010000000011011;
		#400 //4.2340474e+33 * 8.530592e-15 = 3.6118928e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010001011001001111101000110010;
		b = 32'b01000111000001110100010011010110;
		correct = 32'b01011000111100011111101100000100;
		#400 //61465633000.0 * 34628.836 = 2128483200000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000110101100110010001110110;
		b = 32'b00110010011001001111011001101011;
		correct = 32'b10100011101111111011111111010111;
		#400 //-1.5599102e-09 * 1.3327376e-08 = -2.0789509e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101101010000001101010100101111;
		b = 32'b10011010011001110110010000101101;
		correct = 32'b01001000001011100100101111010011;
		#400 //-3.7299278e+27 * -4.7850602e-23 = 178479.3
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110101111000001010111111010000;
		b = 32'b01000010010001111010111111010101;
		correct = 32'b10111000101011110100001011111110;
		#400 //-1.6740469e-06 * 49.92171 = -8.3571285e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101000011011010011111011011111;
		b = 32'b10100010110011001101100001010111;
		correct = 32'b11001011101111011101011010010111;
		#400 //4.4814425e+24 * -5.552337e-18 = -24882478.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000100111101010001010101110110;
		b = 32'b01110111011011100111001001100010;
		correct = 32'b10111100111001000100011101110101;
		#400 //-5.7618932e-36 * 4.8362758e+33 = -0.027866105
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001100111001011001010110001111;
		b = 32'b10011100011100110010101001000001;
		correct = 32'b10101001110110100001001011011100;
		#400 //120368250.0 * -8.0456567e-22 = -9.6844164e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100100100100111110001011010010;
		b = 32'b10010001000001010100010101011100;
		correct = 32'b10110110000110011111100111010001;
		#400 //2.1824124e+22 * -1.0513223e-28 = -2.294419e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001000100010111111011100101010;
		b = 32'b11110010101000000111101111000110;
		correct = 32'b01111011101011110111110001001101;
		#400 //-286649.3 * -6.357406e+30 = 1.8223461e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111001100100100010011111110100;
		b = 32'b00010001010111011101011011100000;
		correct = 32'b11001011011111010100111001010110;
		#400 //-9.486071e+34 * 1.750004e-28 = -16600662.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111011000100100000000110001;
		b = 32'b11001011000100111011011011000111;
		correct = 32'b01000011000000101000110001100110;
		#400 //-1.3485595e-05 * -9680583.0 = 130.54843
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010100011010110010101110101111;
		b = 32'b01100101010100010011001011100000;
		correct = 32'b01111010010000000010110101100110;
		#400 //4040200800000.0 * 6.1744567e+22 = 2.4946045e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111101101001010100101010111;
		b = 32'b10100111100011011000100000111110;
		correct = 32'b10101111110001111100001011010101;
		#400 //92498.68 * -3.9283076e-15 = -3.6336326e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111011111010000100010000010000;
		b = 32'b01110001110000101001011100100111;
		correct = 32'b01101110001100001000110010111000;
		#400 //0.007088192 * 1.9271304e+30 = 1.365987e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001100011010000011101001101010;
		b = 32'b11011111001001101011010111010111;
		correct = 32'b11101100000101110011101011010101;
		#400 //60877224.0 * -1.2012744e+19 = -7.313025e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111101100111110000100100110000;
		b = 32'b00001101011001100110100111101010;
		correct = 32'b01001011100011110010010000001101;
		#400 //2.642437e+37 * 7.100171e-31 = 18761754.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011101011110000011000010010010;
		b = 32'b01111010011011011100101110101101;
		correct = 32'b01011000011001101000101001101101;
		#400 //3.2847637e-21 * 3.0867635e+35 = 1013928830000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111110000101001000111001011100;
		b = 32'b10111101101000010111001010011001;
		correct = 32'b11111100001110110110000000010000;
		#400 //4.936623e+37 * -0.07883186 = -3.8916316e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100011101010001010001111001101;
		b = 32'b11101000000011101010000001110110;
		correct = 32'b01001100001110111110100100100000;
		#400 //-1.8283969e-17 * -2.694144e+24 = 49259650.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101101000100010111010000110100;
		b = 32'b01000001100110001111110111101110;
		correct = 32'b10101111001011011101101010001100;
		#400 //-8.268098e-12 * 19.12399 = -1.5811902e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010100010101100001101001101010;
		b = 32'b10110000001110010100001011110101;
		correct = 32'b00000101000110101111000100010110;
		#400 //-1.0809448e-26 * -6.739776e-10 = 7.285326e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011110010101111100111111101000;
		b = 32'b01011001100110101011010111100110;
		correct = 32'b01111000100000100110110001101001;
		#400 //3.8877258e+18 * 5443393000000000.0 = 2.116242e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000111100101010101001000000110;
		b = 32'b11000010111001110011101110110111;
		correct = 32'b10001011000001101101111111011000;
		#400 //2.2467237e-34 * -115.61663 = -2.5975863e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111000111101011001011000001010;
		b = 32'b00011000011101111010000010001000;
		correct = 32'b00010001111011011000110111000100;
		#400 //0.00011710457 * 3.200505e-24 = 3.7479377e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111001000111110101111111101000;
		b = 32'b00001001000100101001000000111010;
		correct = 32'b10000010101101100111110011111001;
		#400 //-0.0001519915 * 1.7641926e-33 = -2.6814227e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111101110110011011010001111000;
		b = 32'b01010010000101010001010101001110;
		correct = 32'b01010000011111011001000001010000;
		#400 //0.10630125 * 160076890000.0 = 17016373000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101111000000010001011001100000;
		b = 32'b11100011001001000101010001111001;
		correct = 32'b01010010101001011011100111011100;
		#400 //-1.1740431e-10 * -3.031353e+21 = 355893900000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000010110111111111000001100010;
		b = 32'b11111000001110101011101001001010;
		correct = 32'b01111011101000110101011110011101;
		#400 //-111.9695 * -1.514915e+34 = 1.6962428e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110111110101100100011010000101;
		b = 32'b11001001111100110101011101110010;
		correct = 32'b11000010010010111010111000100010;
		#400 //2.5543626e-05 * -1993454.2 = -50.92005
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110100101101001101011101000100;
		b = 32'b01011011011010010001001011011000;
		correct = 32'b11010000101001001010010100111101;
		#400 //-3.368424e-07 * 6.560439e+16 = -22098340000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001010110110101010011111011100;
		b = 32'b11000010011101111111001100101100;
		correct = 32'b00001101110100111100011110101000;
		#400 //-2.1055778e-32 * -61.987473 = 1.30519445e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111110101110101000011110110111;
		b = 32'b00011110011001000100100000011011;
		correct = 32'b11011101101001100101010101101001;
		#400 //-1.2397054e+38 * 1.20851306e-20 = -1.4982002e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000101100010110100001110100110;
		b = 32'b01010111001000001010101111011111;
		correct = 32'b10011101001011101100111110001110;
		#400 //-1.3096347e-35 * 176660040000000.0 = -2.3136012e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100101010100001010111000101111;
		b = 32'b01010111010010000011001011101111;
		correct = 32'b10111101001000110011000110011010;
		#400 //-1.810014e-16 * 220121080000000.0 = -0.039842226
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110001100100001100001011110010;
		b = 32'b00101110001111000101100001010111;
		correct = 32'b01100000010101010000001000111100;
		#400 //1.4336485e+30 * 4.2824713e-11 = 6.1395586e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000011010001001101000010010100;
		b = 32'b00010011010100100110011111011010;
		correct = 32'b10010111001000011100001011110001;
		#400 //-196.81476 * 2.655693e-27 = -5.2267956e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111001100010111000011000100011;
		b = 32'b11011000110110101101001111011100;
		correct = 32'b01010010111011101000011101100011;
		#400 //-0.00026612086 * -1924827700000000.0 = 512236800000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100000111101010100101001011000;
		b = 32'b11100110000011110101101111100101;
		correct = 32'b01000111100010010101110010010100;
		#400 //-4.155381e-19 * -1.6924839e+23 = 70329.16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000101000011011100100001000110;
		b = 32'b01110010110111110011010011100001;
		correct = 32'b00111000011101110011110101111101;
		#400 //6.6665726e-36 * 8.842123e+30 = 5.8946654e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010011100101101111101100110001;
		b = 32'b01110111001000101111010010100001;
		correct = 32'b01001011010000000011011001110111;
		#400 //3.8113017e-27 * 3.305132e+33 = 12596855.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011110100110001000100111011001;
		b = 32'b10000001000100010010100010101010;
		correct = 32'b10100000001011001111110010011101;
		#400 //5.4957775e+18 * -2.666147e-38 = -1.465255e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100010010100001011111101110111;
		b = 32'b11111100000001100101111000010111;
		correct = 32'b11011110110110110010000111100011;
		#400 //2.8290617e-18 * -2.7907046e+36 = -7.8950757e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111111001000111000101100010;
		b = 32'b10001101101111011111111101000010;
		correct = 32'b00000110001010011000101101111101;
		#400 //-2.7232516e-05 * -1.1709475e-30 = 3.1887847e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101110100101001001010110000011;
		b = 32'b10101011111010111001101101101011;
		correct = 32'b01011011000010001011111101110100;
		#400 //-2.2992265e+28 * -1.6740891e-12 = 3.84911e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111000010010000101100100011110;
		b = 32'b11000100011001010101001100100111;
		correct = 32'b01111101001100110111100011001011;
		#400 //-1.625417e+34 * -917.29926 = 1.4909938e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110101001100110001001111001110;
		b = 32'b00010001000110011111110110000100;
		correct = 32'b01000110110101110111000001011010;
		#400 //2.2700753e+32 * 1.2147692e-28 = 27576.176
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110011100000111011011001101000;
		b = 32'b01110100011001011110010110111000;
		correct = 32'b01101000011011001001000010111000;
		#400 //6.1333424e-08 * 7.2857375e+31 = 4.4685923e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101110011110101100011001010011;
		b = 32'b11001010010111000111101011100100;
		correct = 32'b01111001010101111111101011010001;
		#400 //-1.9402753e+28 * -3612345.0 = 7.0089437e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000010100100101100111000111000;
		b = 32'b01000000000100101100110001111010;
		correct = 32'b01000011001010000101110110111100;
		#400 //73.40277 * 2.2937303 = 168.36615
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100110101001011011000110010101;
		b = 32'b01000110000011011000111001100100;
		correct = 32'b11101101001101110011110111110001;
		#400 //-3.9123314e+23 * 9059.598 = -3.544415e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100110111110101010110011000100;
		b = 32'b00101101101100111010011111010111;
		correct = 32'b11010101001011111110101100100110;
		#400 //-5.918893e+23 * 2.042448e-11 = -12089031000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110100100111000110011110110001;
		b = 32'b10011011100100011110100101000001;
		correct = 32'b00010000101100100100101001111011;
		#400 //-2.913271e-07 * -2.4138975e-22 = 7.0323376e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000101000011011100110001000011;
		b = 32'b00000101100111111010100010011010;
		correct = 32'b00001011001100001101111010000010;
		#400 //2268.7664 * 1.5014223e-35 = 3.4063763e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111010100101111101100000000110;
		b = 32'b00001100101110101010010011111101;
		correct = 32'b00000111110111010110100110100010;
		#400 //0.0011584766 * 2.8757136e-31 = 3.331447e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100011110010011011010111111011;
		b = 32'b01000111100100101011111011111101;
		correct = 32'b01101011111001110100000010001011;
		#400 //7.441817e+21 * 75133.98 = 5.5913332e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100010100011010001101110110010;
		b = 32'b10001001111010101010100010010110;
		correct = 32'b00101101000000010101100000111110;
		#400 //-1.3014933e+21 * -5.649199e-33 = 7.352395e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010001101111001111110101111111;
		b = 32'b11110100110010001111001111101110;
		correct = 32'b01000111000101000101101000100000;
		#400 //-2.98174e-28 * -1.27369e+32 = 37978.125
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101001001101001111000100001111;
		b = 32'b00001000111111010100001100101000;
		correct = 32'b00110010101100110000000110110011;
		#400 //1.3671563e+25 * 1.5242672e-33 = 2.0839115e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010110110101111011101000000000;
		b = 32'b10011011011100011101000110100101;
		correct = 32'b00110010110010111100011011000100;
		#400 //-118596930000000.0 * -2.0002793e-22 = 2.3722698e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000101101100110000111100111011;
		b = 32'b01011011000001101111100010100011;
		correct = 32'b00100001001111001100111111000011;
		#400 //1.6838674e-35 * 3.7991026e+16 = 6.397185e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100101110110111010000100001101;
		b = 32'b10000000000110010100110110111110;
		correct = 32'b00100101101011011010101101100110;
		#400 //-1.2964614e+23 * -2.323776e-39 = 3.012686e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110101101010001110001001000001;
		b = 32'b01111101110111011010010011011010;
		correct = 32'b01110100000100100011100000010011;
		#400 //1.2582824e-06 * 3.6826918e+37 = 4.6338663e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011110011110010010010000000001;
		b = 32'b10101101101010111011101100111001;
		correct = 32'b11001100101001110010000101000001;
		#400 //4.4881188e+18 * -1.9523593e-11 = -87624200.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000101101101100011100110000110;
		b = 32'b11100101110011011110100111101000;
		correct = 32'b10101100000100101001001010010000;
		#400 //1.7136329e-35 * -1.2154999e+23 = -2.0829206e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100111101011101000101101111;
		b = 32'b11001001010110001000010000000111;
		correct = 32'b11001110110011111110011101111100;
		#400 //1966.5448 * -886848.44 = -1744027100.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101001110000111100011111011001;
		b = 32'b10011011000100001001111110101000;
		correct = 32'b01000101010111010011010100000111;
		#400 //-2.9585536e+25 * -1.1962989e-22 = 3539.3142
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011010101101101110010100000100;
		b = 32'b01011011000101011011110100000001;
		correct = 32'b01110110010101011111010010100110;
		#400 //2.5740126e+16 * 4.2147584e+16 = 1.0848841e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110100111111101100110010001000;
		b = 32'b10001101110100111011010101111001;
		correct = 32'b00000011010100101011011100110011;
		#400 //-4.7460003e-07 * -1.3047567e-30 = 6.1923756e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100101000110011101100111110101;
		b = 32'b00001011011011011101000001011101;
		correct = 32'b00110001000011101110110000000001;
		#400 //4.5408917e+22 * 4.5801295e-32 = 2.0797872e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011011100111101100111111000001;
		b = 32'b10010111110001001111001010011111;
		correct = 32'b00110011111101000101101100100110;
		#400 //-8.940295e+16 * -1.2727449e-24 = 1.1378715e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001001010011101110101101110000;
		b = 32'b11101010100100110001011011011001;
		correct = 32'b11110100011011011100011101010010;
		#400 //847543.0 * -8.8909995e+25 = -7.5355045e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010111011111001010000101100101;
		b = 32'b10110111110101111101100101000100;
		correct = 32'b01001111110101010000000111110100;
		#400 //-277770110000000.0 * -2.573117e-05 = 7147350000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110001100011110011111010010100;
		b = 32'b10011100101000100000001001110000;
		correct = 32'b01001110101101010100110111101110;
		#400 //-1.4186243e+30 * -1.0720891e-21 = 1520891600.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000110101011111000010010100101;
		b = 32'b11011011111011000011011001011011;
		correct = 32'b11100011001000011111001110001100;
		#400 //22466.322 * -1.3297572e+17 = -2.9874752e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110000100011011110010101000;
		b = 32'b00110011011010010100111001100000;
		correct = 32'b00110010000001001101000101010011;
		#400 //0.14232123 * 5.432082e-08 = 7.731006e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100010011011111001011101000000;
		b = 32'b11101000101110111000101000111001;
		correct = 32'b11001011101011111000010011011001;
		#400 //3.247061e-18 * -7.0850583e+24 = -23005618.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110001011010000101001110101111;
		b = 32'b10110011111110111100001101111100;
		correct = 32'b01100101111001000111101101110101;
		#400 //-1.150427e+30 * -1.1723657e-07 = 1.3487212e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000110111000011010100111101010;
		b = 32'b01010110011110110010110111001011;
		correct = 32'b11011101110111010110100111110110;
		#400 //-28884.957 * 69043524000000.0 = -1.9943192e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010111100110010011010000011001;
		b = 32'b01100000001101000111001110101011;
		correct = 32'b00111000010101111111101110110101;
		#400 //9.900545e-25 * 5.20117e+19 = 5.1494415e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111101010000000001001101111011;
		b = 32'b00101010001100110101011001110011;
		correct = 32'b11101000000001101000111001111100;
		#400 //-1.5957058e+37 * 1.5928387e-13 = -2.541702e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011110110101000101101011111101;
		b = 32'b01100100001000101111111101101111;
		correct = 32'b11000011100001110011010101110111;
		#400 //-2.2484005e-20 * 1.2027114e+22 = -270.4177
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010110010101110001011000101010;
		b = 32'b00000000010100101101110100110010;
		correct = 32'b10010111000010110011110111100011;
		#400 //-59122550000000.0 * 7.60986e-39 = -4.4991434e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110100101101001001101011101111;
		b = 32'b00100010111001001110100001011000;
		correct = 32'b10011000001000010111110111100111;
		#400 //-3.3640342e-07 * 6.2045527e-18 = -2.0872327e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111000110011011001000101101111;
		b = 32'b01111101011000000000010100111010;
		correct = 32'b01110110101100111110001101110100;
		#400 //9.802251e-05 * 1.8610888e+37 = 1.824286e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010101011110001001001111111111;
		b = 32'b10110111000000001000000101010100;
		correct = 32'b01001100111110011000111100100111;
		#400 //-17082158000000.0 * -7.659506e-06 = 130840890.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111100100001011010000100101111;
		b = 32'b00010100100110111110101110000011;
		correct = 32'b01010001101000101100011100001110;
		#400 //5.5507574e+36 * 1.5743893e-26 = 87390536000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110101010011110110110100110001;
		b = 32'b10100110001111101011110000011100;
		correct = 32'b00011100000110101000101101110101;
		#400 //-7.7272404e-07 * -6.617443e-16 = 5.113457e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001110111010111011110111100010;
		b = 32'b01100010110111011000000001000111;
		correct = 32'b11110010010010111111100100001100;
		#400 //-1977545000.0 * 2.0429869e+21 = -4.0400983e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100010110111101011100111010;
		b = 32'b10000011110000100111001101101000;
		correct = 32'b10001000101001101111110000110101;
		#400 //879.3629 * -1.1428791e-36 = -1.0050055e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100001111011110010000010010;
		b = 32'b01110010110110001010110111010001;
		correct = 32'b01110111101000001011100101011101;
		#400 //759.5636 * 8.5835383e+30 = 6.519743e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101110101000110011100000110110;
		b = 32'b00010110001011000100000001010000;
		correct = 32'b01000101010110111010010110001011;
		#400 //2.5257006e+28 * 1.3914343e-25 = 3514.3464
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011011111111110110000110001001;
		b = 32'b00110111101100101100011011011000;
		correct = 32'b01010100001100100101100000101110;
		#400 //1.4376672e+17 * 2.1311847e-05 = 3063934400000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111111011111011000100101000011;
		b = 32'b10100101101000000101100111010110;
		correct = 32'b00100101100111101100111011000011;
		#400 //-0.9903757 * -2.781645e-16 = 2.7548738e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011100010010000111101111101010;
		b = 32'b10010010000010000011000100111100;
		correct = 32'b00101110110101010101000011000110;
		#400 //-2.2572496e+17 * -4.297472e-28 = 9.700467e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001000001100101101100100001001;
		b = 32'b10000000011010011011000000111010;
		correct = 32'b10001001000100111010110001000101;
		#400 //183140.14 * -9.705945e-39 = -1.7775482e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111101011100011011000101001101;
		b = 32'b10010110101110101001101000010001;
		correct = 32'b11010100101100000010110001000111;
		#400 //2.0079034e+37 * -3.014715e-25 = -6053257000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000111000100100111010000010110;
		b = 32'b11100111111010101000110000010100;
		correct = 32'b10101111100001100010111000111111;
		#400 //1.1017934e-34 * -2.2152355e+24 = -2.4407318e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111001010110011001001110110101;
		b = 32'b00010111001010111100001101000111;
		correct = 32'b01010001000100011111101110100010;
		#400 //7.0607767e+34 * 5.5499555e-25 = 39186997000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001100000010110101110100101011;
		b = 32'b10111110001111100101111100110010;
		correct = 32'b10001010110011110100010111110001;
		#400 //1.0736207e-31 * -0.18591002 = -1.9959684e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001111000011110001111101111110;
		b = 32'b00101001010011101111010110001011;
		correct = 32'b00111000111001110110100100111100;
		#400 //2401205800.0 * 4.5954163e-14 = 0.0001103454
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110001111101011001010001010110;
		b = 32'b00011000011111000011010010101011;
		correct = 32'b10001010111100011111000010001011;
		#400 //-7.1473023e-09 * 3.2596827e-24 = -2.3297938e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100101100100110011101101100010;
		b = 32'b00100001001010101101010101001111;
		correct = 32'b10000111010001001000000000111010;
		#400 //-2.5540674e-16 * 5.788055e-19 = -1.4783084e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100110111001111011111100111100;
		b = 32'b01000111111011111110010011101000;
		correct = 32'b10101111010110010010101011000001;
		#400 //-1.6080679e-15 * 122825.81 = -1.9751224e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010010110111101000100011011110;
		b = 32'b01100001110001010011111101000110;
		correct = 32'b10110101001010110111011001010011;
		#400 //-1.404391e-27 * 4.54821e+20 = -6.387465e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011110101101100110101001011001;
		b = 32'b10001101100001010101000100010011;
		correct = 32'b00101100101111011111111000001011;
		#400 //-6.572208e+18 * -8.216276e-31 = 5.3999075e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111101110011010110110000001010;
		b = 32'b10010110000110011011001010011110;
		correct = 32'b10010100011101101010100111001100;
		#400 //0.100303724 * -1.2415603e-25 = -1.2453313e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001010100101110010000001010001;
		b = 32'b10100111000101001101111100110110;
		correct = 32'b00110010001011111100010011101000;
		#400 //-4952104.5 * -2.0660129e-15 = 1.0231112e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111000001011000110100110001011;
		b = 32'b10010011101010111011111001000001;
		correct = 32'b11001100011001110101010101000100;
		#400 //1.3987746e+34 * -4.3354074e-27 = -60642576.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000010110111011001001110101000;
		b = 32'b10101100011001010110110110110110;
		correct = 32'b00101111110001101001010000001011;
		#400 //-110.78839 * -3.260376e-12 = 3.612118e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010001101000000110001011111100;
		b = 32'b01000000100110110001110010011100;
		correct = 32'b11010010110000100101101110110110;
		#400 //-86106930000.0 * 4.8472424 = -417381150000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010110010010011101011101000111;
		b = 32'b10101001111100011100111010011101;
		correct = 32'b10000000101111101010011010010001;
		#400 //1.630458e-25 * -1.07383916e-13 = -1.7508497e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101101100101101100011011101111;
		b = 32'b01101000010001000000100010001001;
		correct = 32'b01010110011001101110101010101100;
		#400 //1.714137e-11 * 3.702965e+24 = 63473896000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110000010011100000000001001111;
		b = 32'b10110000101100100111001001100011;
		correct = 32'b01100001100011111001100001000011;
		#400 //-2.5501714e+29 * -1.2983715e-09 = 3.31107e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110001110001000000001111001100;
		b = 32'b10100101110100010110101010101110;
		correct = 32'b01011000001000000101100011001000;
		#400 //-1.9412369e+30 * -3.632801e-16 = 705212700000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011111011110001111101100000001;
		b = 32'b11010101111100011111011110000100;
		correct = 32'b11110101111010110101010100000111;
		#400 //1.7940935e+19 * -33255672000000.0 = -5.9663785e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001010000010111011110111101001;
		b = 32'b01001010010100110011111001010000;
		correct = 32'b10010100111001101001111100010101;
		#400 //-6.728325e-33 * 3461012.0 = -2.3286812e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110101011110011100000101001101;
		b = 32'b11100111010000001001111000011100;
		correct = 32'b01011101001110111110101100111010;
		#400 //-9.304102e-07 * -9.09611e+23 = 8.463113e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100110101011101111110100011000;
		b = 32'b11000111100100111011110110101001;
		correct = 32'b11101110110010011111100111110010;
		#400 //4.1318026e+23 * -75643.32 = -3.1254326e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101111011001101110010011111110;
		b = 32'b10111100100101010010000000101000;
		correct = 32'b11101100100001101000000001001001;
		#400 //7.1458387e+28 * -0.01820381 = -1.300815e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001110100001000001001101101001;
		b = 32'b01000100111010001001110001111100;
		correct = 32'b11010011111100000000010010100110;
		#400 //-1107932300.0 * 1860.8901 = -2061740300000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010000100011110001111010000101;
		b = 32'b10101010111001000100111110100110;
		correct = 32'b10111011111111110100011101101011;
		#400 //19209136000.0 * -4.0556203e-13 = -0.007790496
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100010100110100110000000100001;
		b = 32'b01010100011100001100111111111111;
		correct = 32'b10110111100100010011011110001100;
		#400 //-4.1843564e-18 * 4137127000000.0 = -1.7311213e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101001000000110010000111101101;
		b = 32'b11101110100001011011010101111111;
		correct = 32'b11011000000010001111101100110000;
		#400 //2.911727e-14 * -2.069046e+28 = -602449700000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101011100001100100011101000101;
		b = 32'b00100001000100111111001101110111;
		correct = 32'b00001101000110110011010101000001;
		#400 //9.541054e-13 * 5.012776e-19 = 4.7827165e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001100011100110001101000110100;
		b = 32'b01100001010001001011110000100111;
		correct = 32'b00101110001110101101001010111100;
		#400 //1.8727924e-31 * 2.2681998e+20 = 4.2478673e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111101011001001001000011101100;
		b = 32'b00010011100000101010111100010111;
		correct = 32'b11010001011010010101101111010111;
		#400 //-1.8988529e+37 * 3.2989266e-27 = -62641762000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001010001101011010110110000101;
		b = 32'b01110100011010110011000011111011;
		correct = 32'b01111111001001101110100100001100;
		#400 //2976609.2 * 7.453511e+31 = 2.218619e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110010001011111000011000010000;
		b = 32'b10010101101101111111101101111100;
		correct = 32'b10001000011111000100101010000110;
		#400 //1.0216823e-08 * -7.4309884e-26 = -7.5921093e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110111000100101000100110001001;
		b = 32'b10001100010101000110100011011010;
		correct = 32'b01000011111100110010101111010100;
		#400 //-2.9721285e+33 * -1.6363439e-31 = 486.3424
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100100100000010100000011001000;
		b = 32'b11100000001111001010101000011000;
		correct = 32'b11000101001111101000001011101000;
		#400 //5.6054576e-17 * -5.437882e+19 = -3048.1816
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100001011110000111011010100110;
		b = 32'b10110100111101100010010111101101;
		correct = 32'b00010110111011101110011011010011;
		#400 //-8.41827e-19 * -4.5848665e-07 = 3.8596644e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101010101111111110101101010101;
		b = 32'b00100111010101010100000101000100;
		correct = 32'b11010010100111111101111110111011;
		#400 //-1.1600808e+26 * 2.9595069e-15 = -343326700000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111100101111111100100011100010;
		b = 32'b00100011011110011001100101010000;
		correct = 32'b01100000101110101111110100111111;
		#400 //7.966425e+36 * 1.3530782e-17 = 1.0779196e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010100000100110110000100010001;
		b = 32'b00101110100010011100011010000101;
		correct = 32'b00000011000111101010001001110111;
		#400 //7.440746e-27 * 6.265303e-11 = 4.6618527e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101111000110110100101010010111;
		b = 32'b01111101111110011100011100110101;
		correct = 32'b11101101100101111000010001100100;
		#400 //-1.4123668e-10 * 4.1501514e+37 = -5.861536e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101001011111100110111000110010;
		b = 32'b11111111111010001100100101111101;
		correct = 32'b11111111111010001100100101111101;
		#400 //-1.9224221e+25 * nan = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100000101101111011111100110001;
		b = 32'b01100100100111000101101110111100;
		correct = 32'b11000101111000000111010010110100;
		#400 //-3.1127926e-19 * 2.3074418e+22 = -7182.588
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101010111101111011101100011100;
		b = 32'b11111110101000010101110001101000;
		correct = 32'b01101010000111000010011000011000;
		#400 //-4.4005847e-13 * -1.0724275e+38 = 4.719308e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010011001101010011111011000000;
		b = 32'b00000001101011000111111000000100;
		correct = 32'b10010101011101000011111011000001;
		#400 //-778441850000.0 * 6.3363645e-38 = -4.9324912e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011101010001110011111011000100;
		b = 32'b10100111000001000111110110100101;
		correct = 32'b11000100110011100011110001001110;
		#400 //8.973205e+17 * -1.8386792e-15 = -1649.8845
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011010110001011001101001110111;
		b = 32'b01011111101111100011111010011101;
		correct = 32'b01111011000100101101100011111001;
		#400 //2.7810203e+16 * 2.7417134e+19 = 7.624761e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110000100001110101001111111010;
		b = 32'b10010011011001011010110110000111;
		correct = 32'b01000100011100101101001110110011;
		#400 //-3.35056e+29 * -2.898942e-27 = 971.3078
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000110110001010011010110101001;
		b = 32'b11101000110011001110101101101010;
		correct = 32'b11110000000111011101110000011101;
		#400 //25242.83 * -7.741643e+24 = -1.9542099e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011011010100111001110001111111;
		b = 32'b01010011100010111100111000111101;
		correct = 32'b11101111011001110010000011100111;
		#400 //-5.956329e+16 * 1200921100000.0 = -7.1530814e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010010111101101010011100101111;
		b = 32'b00001010100111101011010011101000;
		correct = 32'b00011110000110001110100101111100;
		#400 //529683400000.0 * 1.5282896e-32 = 8.0950964e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000010110011110110110100100011;
		b = 32'b01110001100111111110001000010101;
		correct = 32'b11110101000000011000101111111000;
		#400 //-103.71316 * 1.5834059e+30 = -1.6422002e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001000000001001111001001111010;
		b = 32'b10111010101010010101101111000000;
		correct = 32'b01000011001011111110011101110001;
		#400 //-136137.9 * -0.001292102 = 175.90407
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001001001110001110111111011111;
		b = 32'b10110001100001010111100000100110;
		correct = 32'b00111011010000001101011011010101;
		#400 //-757501.94 * -3.8844687e-09 = 0.0029424925
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110001011111010111011010110010;
		b = 32'b01011110100111011111111100101100;
		correct = 32'b01010000100111000110111001110000;
		#400 //3.6883816e-09 * 5.6924334e+18 = 20995867000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000110001101010110100000001100;
		b = 32'b01010100101011001110010101000111;
		correct = 32'b01011011011101010000100011000001;
		#400 //11610.012 * 5940648000000.0 = 6.8970994e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011001001110011001000101101110;
		b = 32'b10101101000101010111100110001000;
		correct = 32'b11000110110110001011001101111011;
		#400 //3264548300000000.0 * -8.496655e-12 = -27737.74
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111100011000111101010010100000;
		b = 32'b11101101100010101111110000001111;
		correct = 32'b11101010011101110110000111100010;
		#400 //0.013905674 * -5.3767064e+27 = -7.476673e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110111010111101001101000000110;
		b = 32'b00011000000100001011110111110001;
		correct = 32'b00001111111110111011011110011001;
		#400 //1.32680925e-05 * 1.870746e-24 = 2.482123e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110100000011010101110001101100;
		b = 32'b00101111101111001001011011010100;
		correct = 32'b00100100010100000100011001010001;
		#400 //1.3165271e-07 * 3.430417e-10 = 4.516237e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001100001111111100110101110101;
		b = 32'b11100010000100110010111101010011;
		correct = 32'b10101110110111001000110011011110;
		#400 //1.4775932e-31 * -6.7877036e+20 = -1.0029465e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101001001010010110010000011000;
		b = 32'b00101110111100011100101011000001;
		correct = 32'b10011000100111111111110101100011;
		#400 //-3.7612356e-14 * 1.09954275e-10 = -4.135639e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111011100100011111001010000110;
		b = 32'b10011011110011000000110111100010;
		correct = 32'b01010111111010001010101001011010;
		#400 //-1.515604e+36 * -3.375794e-22 = 511636700000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010101101000011010000010110000;
		b = 32'b00100100010011100100001110111011;
		correct = 32'b00111010100000100011101000010001;
		#400 //22213940000000.0 * 4.47265e-17 = 0.0009935518
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101000001100000001010100110000;
		b = 32'b11000010101001111110101000000011;
		correct = 32'b10101011011001101111110110001111;
		#400 //9.774557e-15 * -83.957054 = -8.20643e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111011011101000110011000101011;
		b = 32'b01100010100100111101001100111110;
		correct = 32'b11011110100011010010000001010110;
		#400 //-0.0037292342 * 1.3634465e+21 = -5.084611e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100100100101110111011000000011;
		b = 32'b00100110100000101010110010110100;
		correct = 32'b01001011100110101010000000110111;
		#400 //2.2351696e+22 * 9.067373e-16 = 20267118.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101111011111001111101011101011;
		b = 32'b00011110110010100101000110001101;
		correct = 32'b10001110110001111110111010010100;
		#400 //-2.300841e-10 * 2.142131e-20 = -4.928703e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011110001011010111011011001001;
		b = 32'b11000001110000111100011110101011;
		correct = 32'b10100000100001001010100011000110;
		#400 //9.183108e-21 * -24.472494 = -2.2473355e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101000010111011111111001101001;
		b = 32'b10101101101010001010100101011110;
		correct = 32'b10010110100100100100000111010011;
		#400 //1.2323131e-14 * -1.9174603e-11 = -2.3629113e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011111100101111110100110001001;
		b = 32'b11001010111101010111101001100011;
		correct = 32'b11101011000100011010101100100000;
		#400 //2.1892862e+19 * -8043825.5 = -1.7610236e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011100100110011000111000110101;
		b = 32'b11100111100110001010100111000011;
		correct = 32'b11000100101101110010010010000111;
		#400 //1.016145e-21 * -1.4418625e+24 = -1465.1415
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111101000000010010010010111001;
		b = 32'b00111001111001101011111011100000;
		correct = 32'b10110111011010001100111010010001;
		#400 //-0.031529162 * 0.00044011232 = -1.3876373e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011100001001000010011110101110;
		b = 32'b10111010111101001000011100000101;
		correct = 32'b00010111100111001100110001100110;
		#400 //-5.4314333e-22 * -0.0018655962 = 1.0132861e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110101010010001011001110011111;
		b = 32'b10000110000011000001100001010110;
		correct = 32'b00111011110110111010101010011110;
		#400 //-2.5441956e+32 * -2.6348953e-35 = 0.0067036888
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001010011101111001001001110100;
		b = 32'b00001110110110011100100000000110;
		correct = 32'b10011001110100101001110010010101;
		#400 //-4056221.0 * 5.3687246e-30 = -2.1776734e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100100000110001100110010000010;
		b = 32'b01010101011101111000011110001100;
		correct = 32'b01111010000100111011111000111001;
		#400 //1.1274566e+22 * 17010096000000.0 = 1.9178145e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001101100011001110011001101010;
		b = 32'b01011101010011111100011101011110;
		correct = 32'b10101011011001001011100000010101;
		#400 //-8.683636e-31 * 9.357524e+17 = -8.1257337e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010100011111000101110010101010;
		b = 32'b01010100011001010100010110110101;
		correct = 32'b00101001011000100000001110011011;
		#400 //1.27410234e-26 * 3938868000000.0 = 5.0185208e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001110001111001101110100000110;
		b = 32'b01000011011111011101011001111111;
		correct = 32'b00010010001110110100010010101101;
		#400 //2.3279208e-30 * 253.83788 = 5.9091445e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101100001100001000001111010100;
		b = 32'b01010000100100110010000010010010;
		correct = 32'b10111101010010101110010001010000;
		#400 //-2.5084284e-12 * 19747082000.0 = -0.049534142
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010001100100111010100011101110;
		b = 32'b10110111100010001011101100011101;
		correct = 32'b11001001100111011011101101010111;
		#400 //79274295000.0 * -1.6299595e-05 = -1292138.9
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001101010000001100111011010000;
		b = 32'b10100100110001100100001000001100;
		correct = 32'b00110010100101010101000110110011;
		#400 //-202173700.0 * -8.59807e-17 = 1.7383035e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011101010001000111110101001111;
		b = 32'b10101000000101110011110000001000;
		correct = 32'b00000101111010000010011111111010;
		#400 //-2.6005167e-21 * -8.395201e-15 = 2.183186e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011010100111001100101111110110;
		b = 32'b11100111010110001001110101100000;
		correct = 32'b01000010100001001010110001111011;
		#400 //-6.4849604e-23 * -1.0229342e+24 = 66.336876
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100100010100010100001111100110;
		b = 32'b10101011000111110001101100001010;
		correct = 32'b11010000000000100000111101000110;
		#400 //1.5441048e+22 * -5.652567e-13 = -8728156000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000011110011100110010111000000;
		b = 32'b00100101010111111001110000011110;
		correct = 32'b00101001101101000100100010000000;
		#400 //412.79492 * 1.9395061e-16 = 8.0061825e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001011010100001001111111111110;
		b = 32'b00111101001011000000101110101110;
		correct = 32'b10001001000011000011010100000011;
		#400 //-4.0179708e-32 * 0.042003326 = -1.6876813e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110000101110001001010000111001;
		b = 32'b01001000000010111100100111011110;
		correct = 32'b01111001010010011001010000001111;
		#400 //4.5699546e+29 * 143143.47 = 6.5415916e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001100101010111010011110110010;
		b = 32'b11001011100101100110011000110111;
		correct = 32'b11011000110010011011000110011000;
		#400 //89996690.0 * -19713134.0 = -1774116800000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100111110010001010011111011011;
		b = 32'b10110100000001011110000100111101;
		correct = 32'b00011100010100011101111110000000;
		#400 //-5.569314e-15 * -1.2468531e-07 = 6.9441166e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000101111100010110100010100111;
		b = 32'b00111100000001010101111110110001;
		correct = 32'b11000010011110111000101100110111;
		#400 //-7725.0815 * 0.00814049 = -62.885952
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101111110000111101011000111100;
		b = 32'b11010100010111110000010100001001;
		correct = 32'b01000100101010101001101101111000;
		#400 //-3.5622516e-10 * -3831448700000.0 = 1364.8584
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001001001111110100001001010111;
		b = 32'b00010001111111110000111111011100;
		correct = 32'b10011011101111101000111011101110;
		#400 //-783397.44 * 4.024168e-28 = -3.152523e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110011110101010100001110010;
		b = 32'b11110000100100010011110010011001;
		correct = 32'b11101111100011100011010010111110;
		#400 //0.2447832 * -3.5958868e+29 = -8.802127e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100000111110111110001101101000;
		b = 32'b11000000001000010110011011111111;
		correct = 32'b10100001100111101100111101011100;
		#400 //4.267154e-19 * -2.5219114 = -1.0761384e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010100100111011101000011001100;
		b = 32'b10011110101100110110110011111100;
		correct = 32'b10110011110111010011100001011100;
		#400 //5422503000000.0 * -1.8997437e-20 = -1.0301366e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000111011111011000101010001011;
		b = 32'b11101001001100010010110100000010;
		correct = 32'b01110001001011110111100101011101;
		#400 //-64906.543 * -1.3387026e+25 = 8.689055e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111000010100100101111011001001;
		b = 32'b00010100100000010001010010011101;
		correct = 32'b11001101010101000010010101100111;
		#400 //-1.7067263e+34 * 1.3033802e-26 = -222451310.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010100010100110011100101000010;
		b = 32'b10011100010100000010100100101001;
		correct = 32'b10110001001010111100000001111100;
		#400 //3628795000000.0 * -6.8874625e-22 = -2.499319e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010001111101011110010110111110;
		b = 32'b10100001001101010101111100011000;
		correct = 32'b00110011101011100011011011000111;
		#400 //-132015180000.0 * -6.145104e-19 = 8.11247e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101010111111001110011110100100;
		b = 32'b10011000100010110110101001001101;
		correct = 32'b11000100000010011011101011001010;
		#400 //1.528716e+26 * -3.6037994e-24 = -550.9186
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101111000101010110100110110011;
		b = 32'b10101100000000100110010111110101;
		correct = 32'b10011011100110000011011001011101;
		#400 //1.3589023e-10 * -1.8530709e-12 = -2.5181422e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010110001111010010100011010101;
		b = 32'b00011010110111001011011110110011;
		correct = 32'b10110001101000110001011011010011;
		#400 //-51995767000000.0 * 9.128665e-23 = -4.746519e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010011011101010000100100010010;
		b = 32'b00110001111100100000100110100011;
		correct = 32'b00000101111001111010101111001100;
		#400 //3.092782e-27 * 7.0442225e-09 = 2.1786244e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111000011110010001000110010111;
		b = 32'b01101011100100110101001001110001;
		correct = 32'b11100100100011110101010101001111;
		#400 //-5.9382608e-05 * 3.5620283e+26 = -2.1152252e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101010011000100000101011111010;
		b = 32'b10101111101100000000000111001010;
		correct = 32'b11011010100110110110100100100000;
		#400 //6.8317268e+25 * -3.2015485e-10 = -2.1872104e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111010010100010000110101110110;
		b = 32'b10101100010000011000110000100001;
		correct = 32'b01100111000111100000110110010100;
		#400 //-2.7136577e+35 * -2.7504737e-12 = 7.463844e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111000000001101110000000110101;
		b = 32'b10100011011000110101111100100110;
		correct = 32'b00011011111011111001010111100000;
		#400 //-3.21569e-05 * -1.2325843e-17 = 3.9636088e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000110001100101000110001100010;
		b = 32'b00100111110111000000101101110100;
		correct = 32'b10101110100110010111100010100001;
		#400 //-11427.096 * 6.1074684e-15 = -6.9790625e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101110111011001100010001010011;
		b = 32'b00010011111011001110111011011000;
		correct = 32'b00000011010110110010000111100011;
		#400 //1.0766912e-10 * 5.9810294e-27 = 6.4397216e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111110011001000010110100101110;
		b = 32'b01000101101101000100000100110101;
		correct = 32'b11000100101000001010100111100011;
		#400 //-0.2228286 * 5768.151 = -1285.309
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111001000110110000000110101100;
		b = 32'b10100010111001010100000010000001;
		correct = 32'b00011100100010101100111110001101;
		#400 //-0.00014782575 * -6.213887e-18 = 9.185725e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100000000111101110010110110001;
		b = 32'b01000110110011110000000111101110;
		correct = 32'b00100111100000000111110011101101;
		#400 //1.3459119e-19 * 26496.965 = 3.566258e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100000011001011011100011100111;
		b = 32'b01001011100001011110000000001111;
		correct = 32'b10101100011100000100010000111111;
		#400 //-1.9458234e-19 * 17547294.0 = -3.4143936e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101111110111110101111111001001;
		b = 32'b10000000101010001001111111011110;
		correct = 32'b00110001000100110010001001011010;
		#400 //-1.3826191e+29 * -1.5485713e-38 = 2.1410842e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001010111100100000011010001001;
		b = 32'b11011110100000100101000100110001;
		correct = 32'b01101001111101100110100000101000;
		#400 //-7930692.5 * -4.6951703e+18 = 3.7235952e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100001110010110000001010001000;
		b = 32'b11010100110110001001101110100000;
		correct = 32'b01110111001010111100010110001100;
		#400 //-4.6810893e+20 * -7442591000000.0 = 3.4839433e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000101000111111101000101010110;
		b = 32'b11011011110111011111100001100100;
		correct = 32'b00100001100010101001001011001000;
		#400 //-7.514593e-36 * -1.2495816e+17 = 9.390096e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001100110110010001111110100001;
		b = 32'b01101011101111110010101001101100;
		correct = 32'b10111001001000100010001010010100;
		#400 //-3.345318e-31 * 4.6221033e+26 = -0.00015462405
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010100000001111111010010100100;
		b = 32'b11100000110111010001111011100011;
		correct = 32'b01110101011010101101110100110010;
		#400 //-2335700000000.0 * -1.2746738e+20 = 2.9772555e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010111100001010010010111010001;
		b = 32'b00100110101100111011001111100110;
		correct = 32'b10111110101110101110111000000100;
		#400 //-292794930000000.0 * 1.2469382e-15 = -0.36509717
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110001000001010110100100010101;
		b = 32'b01011011001011000000101110001100;
		correct = 32'b01001100101100110101000100111101;
		#400 //1.941378e-09 * 4.842639e+16 = 94013930.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100101110110011001101110000111;
		b = 32'b10111001111110010111110011101111;
		correct = 32'b11100000010101000001001001111001;
		#400 //1.2845281e+23 * -0.00047586064 = -6.112564e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000000110111111010000101100100;
		b = 32'b10101000111011110001100110101011;
		correct = 32'b10101010010100001101111000011000;
		#400 //6.988451 * -2.6545462e-14 = -1.8551165e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010000000111111010000001101110;
		b = 32'b01001110000000100100101100110000;
		correct = 32'b01011110101000100111110010110100;
		#400 //10712365000.0 * 546491400.0 = 5.8542155e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001010000101101110011010100111;
		b = 32'b00111000011111010101101000111010;
		correct = 32'b01000011000101010101011100100010;
		#400 //2472361.8 * 6.040393e-05 = 149.34036
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010010101010011101111110011011;
		b = 32'b01010111101000101011010110100011;
		correct = 32'b01101010110101111111000000001111;
		#400 //364800480000.0 * 357802000000000.0 = 1.3052635e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011110101110010011000010000001;
		b = 32'b10110011010001110100101001100010;
		correct = 32'b00010010100100000010101010000011;
		#400 //-1.9607698e-20 * -4.640095e-08 = 9.098158e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101001010000111001010001101010;
		b = 32'b01110100010001101100111010001000;
		correct = 32'b11011110000101111110001010010011;
		#400 //-4.3427427e-14 * 6.300438e+31 = -2.736118e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111011110100110110011101001010;
		b = 32'b01110101000110111101000110000110;
		correct = 32'b11110001100000001010110010010000;
		#400 //-0.006451522 * 1.9752335e+32 = -1.2743263e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010101110010100011110110001001;
		b = 32'b10101010011010100001010100010000;
		correct = 32'b11000000101110001110110011100011;
		#400 //27795705000000.0 * -2.0790683e-13 = -5.778917
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101010111100111110011101011011;
		b = 32'b11000011110000101101101011100000;
		correct = 32'b10101111001110011010010111011011;
		#400 //4.3326006e-13 * -389.70996 = -1.6884576e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001010011100001111011111011001;
		b = 32'b00111011110100111001100011111100;
		correct = 32'b11000110110001110010110001001000;
		#400 //-3948022.2 * 0.006457446 = -25494.14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111101111101100111001010001010;
		b = 32'b00110010101110110110001001110010;
		correct = 32'b00110001001101000110010001110000;
		#400 //0.12033565 * 2.1814433e-08 = 2.625054e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101000111010000001110000000011;
		b = 32'b01000001001101010101110111110010;
		correct = 32'b11101010101001000111000011111100;
		#400 //-8.768846e+24 * 11.335436 = -9.939869e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010000101111010110100011011111;
		b = 32'b10011000010001000010001110011011;
		correct = 32'b10101001100100010001111010100011;
		#400 //25422133000.0 * -2.5350382e-24 = -6.444608e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101000010111010000000011001011;
		b = 32'b11001000110101111011000110011100;
		correct = 32'b11110001101110100011010011111111;
		#400 //4.1746305e+24 * -441740.88 = -1.844105e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100100001001110011000000011110;
		b = 32'b00100110010111110110111011000110;
		correct = 32'b00001011000100011110101101000010;
		#400 //3.625311e-17 * 7.7518793e-16 = 2.8102973e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111001101101101011100010110110;
		b = 32'b10101011011001000101010011100111;
		correct = 32'b01100101101000101111100100011100;
		#400 //-1.1859305e+35 * -8.11197e-13 = 9.620233e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001110110000100001111001100101;
		b = 32'b11000111000101111011111000111111;
		correct = 32'b11010110011001100010000001100000;
		#400 //1628385900.0 * -38846.246 = -63256680000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111010100101011011010011111;
		b = 32'b00000001100000100011100000101010;
		correct = 32'b00001001010101100101110111101111;
		#400 //53942.62 * 4.783505e-38 = 2.580348e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101010010101010000100010101110;
		b = 32'b00100010101011100001111000010001;
		correct = 32'b01001101100100001110010011101011;
		#400 //6.4385547e+25 * 4.719463e-18 = 303865180.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100010001000010000001101010010;
		b = 32'b11111000000100101000101111011101;
		correct = 32'b11011010101110000101011110111001;
		#400 //2.1821326e-18 * -1.1889252e+34 = -2.5943924e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000010101001101011000110011111;
		b = 32'b11110100001010010110000011100010;
		correct = 32'b11110111010111001001010010101111;
		#400 //83.34692 * -5.3678173e+31 = -4.47391e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100100100010011111101110001110;
		b = 32'b00110001000100011110001100011001;
		correct = 32'b01010110000111010100001111000110;
		#400 //2.0362643e+22 * 2.1229367e-09 = 43228603000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101010100110101010111100110101;
		b = 32'b00110010000001101100001000011111;
		correct = 32'b00011101001000101101101000000010;
		#400 //2.747747e-13 * 7.843965e-09 = 2.1553229e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101011010100101100011011100100;
		b = 32'b11010000101111110010110001010101;
		correct = 32'b00111100100111010110011011100100;
		#400 //-7.4883003e-13 * -25658829000.0 = 0.019214101
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010000101011100001101110111011;
		b = 32'b00000001111110101111110111010000;
		correct = 32'b00010011001010101011001110110011;
		#400 //23368423000.0 * 9.21997e-38 = 2.1545615e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000001001011000111000111111100;
		b = 32'b11111000101110001110011010111000;
		correct = 32'b11111010011110010001101010101111;
		#400 //10.777828 * -3.0001942e+34 = -3.2335578e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101110111100110101110100110110;
		b = 32'b10011100000101110000101001011110;
		correct = 32'b00001011100011111001010111010110;
		#400 //-1.1066918e-10 * -4.997511e-22 = 5.5307044e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110111110110000110000010001110;
		b = 32'b10101010100000000010011101111010;
		correct = 32'b10100010110110001010001101001010;
		#400 //2.5794168e-05 * -2.276476e-13 = -5.8719806e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101001000100010100101010111100;
		b = 32'b11100110101001100111100001010100;
		correct = 32'b11010000001111001111010110000001;
		#400 //3.226129e-14 * -3.9306625e+23 = -12680824000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110001101101001101001100001101;
		b = 32'b11100110010100111100110001000001;
		correct = 32'b01011000100101011001101000111010;
		#400 //-5.262683e-09 * -2.5004679e+23 = 1315917000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000110011011010000110001001010;
		b = 32'b01001110101011011010010101111111;
		correct = 32'b10010101101000001100101010001101;
		#400 //-4.4583774e-35 * 1456652200.0 = -6.4943054e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100011100010110001010010110011;
		b = 32'b01010111000101001111011101110100;
		correct = 32'b01111011001000011101110011001111;
		#400 //5.131178e+21 * 163790520000000.0 = 8.404383e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111101110101011010011011001001;
		b = 32'b11101010101111110000010000101101;
		correct = 32'b11101001000111110110101011101100;
		#400 //0.10432202 * -1.1546228e+26 = -1.2045258e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001101111001001010110111001000;
		b = 32'b00111010000011110001100111010110;
		correct = 32'b11001000011111111010100001001110;
		#400 //-479574270.0 * 0.0005458867 = -261793.22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110010100111111001101111001111;
		b = 32'b11101100100010110001011111010110;
		correct = 32'b11011111101011010111000011101100;
		#400 //1.858089e-08 * -1.345226e+27 = -2.4995497e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000010010001001111100101010011;
		b = 32'b11100010010000011001000010101100;
		correct = 32'b00100101000101001110111101001000;
		#400 //-1.4471358e-37 * -8.926616e+20 = 1.2918025e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101100011011101111000101100010;
		b = 32'b10010100011011001000000111000101;
		correct = 32'b00000001010111001011111110100110;
		#400 //-3.3955829e-12 * -1.1940548e-26 = 4.054512e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100110000110110010011010111111;
		b = 32'b00011110110010111100101100010000;
		correct = 32'b00000101011101110000010110010110;
		#400 //5.382894e-16 * 2.1577446e-20 = 1.161491e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001000101100001000011110101100;
		b = 32'b01100111001111100010110111110111;
		correct = 32'b11110000100000110010010001100100;
		#400 //-361533.38 * 8.980975e+23 = -3.2469224e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001101111111110010011101110101;
		b = 32'b10010111100001101111000001110101;
		correct = 32'b00100110000001100111111001010001;
		#400 //-535097000.0 * -8.720247e-25 = 4.666178e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010011010101110011101001101010;
		b = 32'b01100010000000101011000000100010;
		correct = 32'b11110101110110111011111101111101;
		#400 //-924398000000.0 * 6.026921e+20 = -5.5712737e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011011000000010000001011010011;
		b = 32'b11101000101110110111100010100000;
		correct = 32'b11000100001111001111001110110100;
		#400 //1.0671542e-22 * -7.0824614e+24 = -755.80786
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010110000111110011001100000010;
		b = 32'b11000001111001000010011010111000;
		correct = 32'b00011000100011011110000110000010;
		#400 //-1.2860013e-25 * -28.518906 = 3.667535e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100010011100101001000001010010;
		b = 32'b01011111111010000100011101111000;
		correct = 32'b11000010110111000001011010000010;
		#400 //-3.2873518e-18 * 3.3474957e+19 = -110.04396
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110101101101111010100011111001;
		b = 32'b01010111111111101000100100010110;
		correct = 32'b01001110001101101001110000000000;
		#400 //1.368374e-06 * 559729470000000.0 = 765919200.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000101001111001100010010010010;
		b = 32'b11111010110010100100100100110001;
		correct = 32'b11000000100101010010100100010011;
		#400 //8.875822e-36 * -5.2516423e+35 = -4.661264
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110100011110011110001010000100;
		b = 32'b10101111000010001111011010101111;
		correct = 32'b00100100000001011011000100100001;
		#400 //-2.3272338e-07 * -1.2456768e-10 = 2.8989812e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101001011101000100101110011000;
		b = 32'b01001101100110000011101110101110;
		correct = 32'b00110111100100010100010111010110;
		#400 //5.424445e-14 * 319256000.0 = 1.7317867e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000110011100100111010001100111;
		b = 32'b01100010111000000100100110111010;
		correct = 32'b11101001110101000110101110101101;
		#400 //-15517.101 * 2.0686916e+21 = -3.2100095e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100001110001110101100110010110;
		b = 32'b01110110001011010001000011110100;
		correct = 32'b01011000100001101100010010111110;
		#400 //1.3508478e-18 * 8.7755e+32 = 1185436500000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011100101100101000001000101110;
		b = 32'b00110101001001001111001100011010;
		correct = 32'b10010010011001100000100111010010;
		#400 //-1.1812703e-21 * 6.144852e-07 = -7.258731e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001000001110111110111001111001;
		b = 32'b10011100111101001100011110111100;
		correct = 32'b00100101101100111011000111101100;
		#400 //-192441.89 * -1.6198196e-21 = 3.1172115e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101101101000001110110100100001;
		b = 32'b00010010100000101101010100001001;
		correct = 32'b10000000101001000111110010101011;
		#400 //-1.82952e-11 * 8.256671e-28 = -1.5105744e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011110110100111100111110110111;
		b = 32'b10111011111001101010011100000011;
		correct = 32'b01011011001111101101011011001101;
		#400 //-7.6313094e+18 * -0.0070389523 = 5.371642e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111000000110011110111011111010;
		b = 32'b11000010100011111100011110000101;
		correct = 32'b00111011001011001110100011101101;
		#400 //-3.6700607e-05 * -71.88969 = 0.0026383952
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001111000001001000010110010101;
		b = 32'b01100000000010010001111100110110;
		correct = 32'b11101111100011011111011101001010;
		#400 //-2223347000.0 * 3.95227e+19 = -8.787268e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111011101101001000001111001;
		b = 32'b01011101000111000011001100100101;
		correct = 32'b01100101000101100111000101001100;
		#400 //63120.473 * 7.034613e+17 = 4.440281e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110101011101110100010000100001;
		b = 32'b00111010100100111100111010010100;
		correct = 32'b00110000100011101100001110100111;
		#400 //9.211381e-07 * 0.0011276775 = 1.0387468e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001010010000110001000000010110;
		b = 32'b10101100000101100011011110010000;
		correct = 32'b00110110111001001110101110000110;
		#400 //-3195909.5 * -2.1347125e-12 = 6.822348e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110110101000011111100000000101;
		b = 32'b00010011111101010000011100001101;
		correct = 32'b01001011000110110000011011010011;
		#400 //1.642559e+33 * 6.1853648e-27 = 10159827.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111101010011001111101111100111;
		b = 32'b00001011001100101011010110011001;
		correct = 32'b10001001000011110001100010001111;
		#400 //-0.05004492 * 3.4418172e-32 = -1.7224546e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011100111010101100110110100011;
		b = 32'b10100011111111110101011011011110;
		correct = 32'b00000001011010100011001010000010;
		#400 //-1.5537977e-21 * -2.7683945e-17 = 4.301525e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001111110100000011111001111011;
		b = 32'b10000010110111010011111001110100;
		correct = 32'b00010011001100111111100010111110;
		#400 //-6987511300.0 * -3.2508878e-37 = 2.2715616e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000110000001011110110101011110;
		b = 32'b00100111011100111100011101100111;
		correct = 32'b10101101111111110001000101000011;
		#400 //-8571.342 * 3.383112e-15 = -2.899781e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000001011110100010101001010101;
		b = 32'b01110010110001010000101101011011;
		correct = 32'b10110100110000001000110110101100;
		#400 //-4.594812e-38 * 7.805731e+30 = -3.5865867e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101000011111111000000001010110;
		b = 32'b00100110110000101101100111000011;
		correct = 32'b10001111110000100111100010011000;
		#400 //-1.4183172e-14 * 1.3520479e-15 = -1.9176328e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011110110110001001011110101110;
		b = 32'b01011110111011011010101111100110;
		correct = 32'b11111110010010010001010111011100;
		#400 //-7.803567e+18 * 8.5630174e+18 = -6.682208e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100110011110110010100011101010;
		b = 32'b01001000001000011111110101100001;
		correct = 32'b11101111000111101110110101010010;
		#400 //-2.9651718e+23 * 165877.52 = -4.9185534e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100101000111010110101001011011;
		b = 32'b11110010100100011010100110010101;
		correct = 32'b01011000001100110010001100001001;
		#400 //-1.3653614e-16 * -5.7702833e+30 = 787852200000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110111010101110101101000101;
		b = 32'b00111110000100111111000011110010;
		correct = 32'b10110101100001111100001000110011;
		#400 //-7.0011324e-06 * 0.14447382 = -1.0114803e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111110111101011110010000100;
		b = 32'b11010001001110100111100000100000;
		correct = 32'b11011001101000100011110101111100;
		#400 //114041.03 * -50054955000.0 = -5708318600000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110101101010010011000110000;
		b = 32'b11101101000110000110010000011011;
		correct = 32'b01100100010101111010101100000101;
		#400 //-5.398666e-06 * -2.9476713e+27 = 1.5913493e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000011001000011011101001101101;
		b = 32'b11110100111000011000100001110010;
		correct = 32'b11111000100011100111101100001101;
		#400 //161.72823 * -1.4294851e+32 = -2.311881e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100101101001110000000101011011;
		b = 32'b01010001101010110000000000001000;
		correct = 32'b10110111110111110001101111011010;
		#400 //-2.89708e-16 * 91804990000.0 = -2.6596641e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000101111100101100011101111010;
		b = 32'b01011101100011011110010100100000;
		correct = 32'b10100100000001101001000100101001;
		#400 //-2.2830847e-35 * 1.2780767e+18 = -2.9179574e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110110000100110001011100110110;
		b = 32'b01110100001111000010000001111100;
		correct = 32'b01101010110110000010111101101100;
		#400 //2.1918217e-06 * 5.961979e+31 = 1.3067596e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111000001111000110000100111110;
		b = 32'b00100110001001100101110010001110;
		correct = 32'b10011110111101001101011001010011;
		#400 //-4.4913257e-05 * 5.7718254e-16 = -2.5923147e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100011101010100000011010010011;
		b = 32'b00110110010100100001011010001110;
		correct = 32'b01011010100010111000100001011111;
		#400 //6.2728404e+21 * 3.1305567e-06 = 1.9637482e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001000111000010001110001010100;
		b = 32'b11001001000100100011111101000111;
		correct = 32'b10010010100000001001100111001100;
		#400 //1.3548355e-33 * -599028.44 = -8.11585e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110110001011101001100111101010;
		b = 32'b00001011001110100010101100111001;
		correct = 32'b00000001111111011111001010011101;
		#400 //2.601761e-06 * 3.5854814e-32 = 9.3285655e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110001100011011101000011110001;
		b = 32'b10100011010111011101010001111110;
		correct = 32'b11010101011101011100011000101110;
		#400 //1.4044794e+30 * -1.2025431e-17 = -16889470000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010101011110101111011000101010;
		b = 32'b00001000011110100110000010110101;
		correct = 32'b00011110011101010111001100110011;
		#400 //17245948000000.0 * 7.5345317e-34 = 1.2994015e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100000111111011000110111010000;
		b = 32'b00110100000001010111110101001010;
		correct = 32'b11010101100001000011011011000101;
		#400 //-1.461639e+20 * 1.243217e-07 = -18171346000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011001001110011010111010100000;
		b = 32'b01111111111101011100110101001001;
		correct = 32'b01111111111101011100110101001001;
		#400 //-3266554600000000.0 * nan = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110100111000100110011011011001;
		b = 32'b00011001001011100010101110011100;
		correct = 32'b01001110100110100000100001111001;
		#400 //1.4349916e+32 * 9.004396e-24 = 1292123300.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011000100010001101110111101011;
		b = 32'b11001101111110101110101001010110;
		correct = 32'b00100111000001100010011000000000;
		#400 //-3.5379256e-24 * -526207680.0 = 1.8616836e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101110010101010000110010011101;
		b = 32'b10111110000100111110110100100011;
		correct = 32'b11101100111101100011011100110000;
		#400 //1.6483889e+28 * -0.14445929 = -2.381251e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000001111111111010011001001100;
		b = 32'b11011001010111110000011110011011;
		correct = 32'b01011011110111101011100101110101;
		#400 //-31.9562 * -3923580000000000.0 = 1.2538271e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110101011001010011010001011010;
		b = 32'b10011000010001111111110100100010;
		correct = 32'b00001110001100110000111001010101;
		#400 //-8.538533e-07 * -2.5847947e-24 = 2.2070354e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011010101000101101011001010110;
		b = 32'b01010001100001100000011100110010;
		correct = 32'b10101100101010101000000110001001;
		#400 //-6.734791e-23 * 71955790000.0 = -4.846072e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010110101000011001100010100110;
		b = 32'b00101001111011000111111111011101;
		correct = 32'b01000001000101010100100101101111;
		#400 //88838500000000.0 * 1.0502686e-13 = 9.330428
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111001100101100011110011111100;
		b = 32'b11000000000011001110001100000011;
		correct = 32'b11111010001001010101110100100111;
		#400 //9.751018e+34 * -2.2013557 = -2.1465458e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111001001101101011101011001011;
		b = 32'b00001011000101001000001010110111;
		correct = 32'b01000100110101000000001010010110;
		#400 //5.9299165e+34 * 2.8602102e-32 = 1696.0808
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101111001011011011110111010011;
		b = 32'b01111100110100101000101000011000;
		correct = 32'b11101100100011101110001101110000;
		#400 //-1.5801697e-10 * 8.745466e+36 = -1.3819321e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001001001011100011001110111111;
		b = 32'b10010101100000100110000110000000;
		correct = 32'b00011111001100010111000100111111;
		#400 //-713531.94 * -5.266041e-26 = 3.7574883e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001101010000111010010110001100;
		b = 32'b01010100111110110100010001000110;
		correct = 32'b01100010110000000000011101111110;
		#400 //205150400.0 * 8633458000000.0 = 1.7711574e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110011101010000111011110000001;
		b = 32'b00100101011100011111001110100011;
		correct = 32'b01011001100111110011100011010101;
		#400 //2.6694632e+31 * 2.0985965e-16 = 5602126000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101100100000110111000000101111;
		b = 32'b11010000110111111110011101001110;
		correct = 32'b00111101111001011110101011110110;
		#400 //-3.735699e-12 * -30051824000.0 = 0.11226456
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100010110101001100110110001001;
		b = 32'b10110110011101000100100110000010;
		correct = 32'b10011001110010110001000100000001;
		#400 //5.7680334e-18 * -3.640162e-06 = -2.0996576e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010010011001010111000100101100;
		b = 32'b00111000111100010010001011101111;
		correct = 32'b00001011110110000001111011011010;
		#400 //7.2399154e-28 * 0.000114982824 = 8.3246594e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100111001100001011011111001011;
		b = 32'b10010100111110010111010000111011;
		correct = 32'b10111100101011000011001100000000;
		#400 //8.345269e+23 * -2.518842e-26 = -0.021020412
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100010101010001111000001110110;
		b = 32'b01100100110000001100010000111110;
		correct = 32'b01000111111111100110101110110011;
		#400 //4.579109e-18 * 2.8447325e+22 = 130263.4
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100100010000001010110110111100;
		b = 32'b00110011100100110000001111111100;
		correct = 32'b00011000010111010100110110000101;
		#400 //4.1780522e-17 * 6.845946e-08 = 2.8602718e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010100100110011010010110100110;
		b = 32'b01011101101111111001000001011000;
		correct = 32'b00110010111001011111001001110010;
		#400 //1.5514389e-26 * 1.7254537e+18 = 2.676936e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111001001001001000010011110111;
		b = 32'b00110000100111110111111110101111;
		correct = 32'b01101010010011010000000101001000;
		#400 //5.3389596e+34 * 1.1605062e-09 = 6.195896e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110000111111011010101111000011;
		b = 32'b10110101011001110101000111000100;
		correct = 32'b01100110111001010011011100000011;
		#400 //-6.2805884e+29 * -8.617319e-07 = 5.4121836e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111101000111010001001000011100;
		b = 32'b00111010000111010010110001000000;
		correct = 32'b01110111110000001101111010000011;
		#400 //1.3048927e+37 * 0.00059956685 = 7.8237037e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000100111100011111100011001000;
		b = 32'b10000010001001101111111000001011;
		correct = 32'b00000111100111011101011101110001;
		#400 //-1935.7744 * -1.2268661e-37 = 2.374936e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011101100001101100000000110101;
		b = 32'b11111111111011110000011011101110;
		correct = 32'b11111111111011110000011011101110;
		#400 //1.2137274e+18 * nan = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001111111001110111001000001011;
		b = 32'b10011101010111011100001001111011;
		correct = 32'b10101101110010000111110101000111;
		#400 //7766021600.0 * -2.934965e-21 = -2.2793002e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100100100111010110101111000110;
		b = 32'b10000011011111000111111101101100;
		correct = 32'b00101000100110110100010001110010;
		#400 //-2.3231238e+22 * -7.4202417e-37 = 1.723814e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101110101111011100010000011011;
		b = 32'b10010111111111100110000110100010;
		correct = 32'b11000111001111001001000011110010;
		#400 //2.9364872e+28 * -1.6439011e-24 = -48272.945
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011011001110110000010110100011;
		b = 32'b00011111011010011100011001110111;
		correct = 32'b00111011001010101100100100011111;
		#400 //5.264202e+16 * 4.9503835e-20 = 0.002605982
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111110011010010111011010100001;
		b = 32'b00011001111001001010111001101011;
		correct = 32'b10011000110100001000110010111000;
		#400 //-0.2279916 * 2.3645094e-23 = -5.390883e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100010010100010000000001110000;
		b = 32'b00101110000000100111101010001011;
		correct = 32'b11010000110101010000110010001001;
		#400 //-9.6385026e+20 * 2.9667418e-11 = -28594948000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111101010111010010010101110101;
		b = 32'b10101001111011010111110100110000;
		correct = 32'b00100111110011010010011111010010;
		#400 //-0.0539908 * -1.0546631e-13 = 5.6942103e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000011110000011011100000010000;
		b = 32'b01001010010010010001101001111010;
		correct = 32'b00001110100110000010110110001110;
		#400 //1.1385779e-36 * 3294878.5 = 3.751476e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110101000111100011111000001111;
		b = 32'b11110101011111010101001101101001;
		correct = 32'b01101011000111001001011011100100;
		#400 //-5.8949894e-07 * -3.2112863e+32 = 1.8930499e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101010101110001101000110101110;
		b = 32'b11110000011110011100100000100100;
		correct = 32'b11011011101101000101010001110000;
		#400 //3.283046e-13 * -3.0921489e+29 = -1.0151667e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101000011100000111110001100011;
		b = 32'b10111010110000110010101010110011;
		correct = 32'b11100011101101110101011011011100;
		#400 //4.54265e+24 * -0.0014890045 = -6.764026e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111001001111010000001001001110;
		b = 32'b00100010010110010011010111111111;
		correct = 32'b00011100001000000101111011010010;
		#400 //0.00018025303 * 2.943757e-18 = 5.306211e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101011111100011101000000010001;
		b = 32'b10100000010101100010000011101111;
		correct = 32'b01001100110010100100001100001010;
		#400 //-5.8466738e+26 * -1.8137402e-19 = 106043470.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101000011010001110100110110110;
		b = 32'b00011101100100011101110000000101;
		correct = 32'b10000110100001001011010010001101;
		#400 //-1.2929265e-14 * 3.8608675e-21 = -4.9918177e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101000000101001000011111111011;
		b = 32'b11011110010000000010010101110001;
		correct = 32'b11000110110111101111011101101011;
		#400 //8.2451364e-15 * -3.4613992e+18 = -28539.709
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001001111100111101110010111110;
		b = 32'b01101000011110011101100001000011;
		correct = 32'b11110010111011011111111110110111;
		#400 //-1997719.8 * 4.7194343e+24 = -9.428107e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110010110000011100001010111110;
		b = 32'b01000111010111111010001000111011;
		correct = 32'b00111010101010010100001101101101;
		#400 //2.2556716e-08 * 57250.23 = 0.0012913771
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000010010001011110101110010010;
		b = 32'b00011001011110111111101101101010;
		correct = 32'b10011100010000101101000001011000;
		#400 //-49.48005 * 1.30271685e-23 = -6.4458494e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001001000100100110100001110100;
		b = 32'b10001000101100011101010110100111;
		correct = 32'b00010010010010110110100011010001;
		#400 //-599687.25 * -1.0703029e-33 = 6.41847e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000110110010011001110000000010;
		b = 32'b11011011101001100110010110100110;
		correct = 32'b10100011000000110000101100110111;
		#400 //7.583703e-35 * -9.367322e+16 = -7.103899e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100111100011101000011001111100;
		b = 32'b00001100000001111010111111011100;
		correct = 32'b10110100000101110001010110101000;
		#400 //-1.3461137e+24 * 1.0452942e-31 = -1.407085e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011101001110010010101111110010;
		b = 32'b11111111010100111010110001110001;
		correct = 32'b01011101000110010001101111110100;
		#400 //-2.4507265e-21 * -2.8136247e+38 = 6.895425e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110111100110110111110000111110;
		b = 32'b11011001000111100111010101001100;
		correct = 32'b11010001010000000111101111011000;
		#400 //1.8535295e-05 * -2787626000000000.0 = -51669467000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111110000110010101100100111100;
		b = 32'b11111100110110111001101001101010;
		correct = 32'b01111011100000111000101111010110;
		#400 //-0.14975446 * -9.121959e+36 = 1.3660542e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010011001000110001110010111;
		b = 32'b01001010101000100001011011000000;
		correct = 32'b11000101100100001001101101010001;
		#400 //-0.000871235 * 5311328.0 = -4627.4146
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011001110101110110101110100001;
		b = 32'b01100110100000100101110100001101;
		correct = 32'b01000000110110110110010111101010;
		#400 //2.227395e-23 * 3.0781206e+23 = 6.8561907
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010110110101101010011000100101;
		b = 32'b10010000100100011010011010111101;
		correct = 32'b10100111111101000011111111010010;
		#400 //118004540000000.0 * -5.7449317e-29 = -6.77928e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011111110010010010011100001110;
		b = 32'b00010001110000111001111101001110;
		correct = 32'b00110010000110011011010111101100;
		#400 //2.8989139e+19 * 3.0863754e-28 = 8.947136e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011111100001011111111011110001;
		b = 32'b11001000010011100010101011000110;
		correct = 32'b10101000010101111101001100010011;
		#400 //5.6749456e-20 * -211115.1 = -1.1980667e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010010100100110001010000100001;
		b = 32'b01011011111101010110001110110111;
		correct = 32'b00101111000011001111101110001110;
		#400 //9.281966e-28 * 1.3814201e+17 = 1.2822296e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100111010010101001000010111110;
		b = 32'b01001000111011001000111010010010;
		correct = 32'b11110000101110110010111000111111;
		#400 //-9.5658805e+23 * 484468.56 = -4.6343684e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010111010001110110110101100011;
		b = 32'b10111100100101010110100011111110;
		correct = 32'b10010100011010001100100011101010;
		#400 //6.4438433e-25 * -0.01823854 = -1.175263e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110111101010000100110100110;
		b = 32'b01000100101011000011001010110011;
		correct = 32'b10111100001001001101001100000011;
		#400 //-7.302692e-06 * 1377.5844 = -0.010060075
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111001101001111110100010111000;
		b = 32'b00101010101010111000100000010011;
		correct = 32'b00100100111000010000001101100110;
		#400 //0.0003202611 * 3.0470122e-13 = 9.758395e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010110010010101011001101110001;
		b = 32'b10101110000000101100000001000001;
		correct = 32'b10000100110011110000111010110011;
		#400 //1.6374052e-25 * -2.9729334e-11 = -4.8678965e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000001111011111100110110110010;
		b = 32'b11010011010111111010001001100000;
		correct = 32'b10010101110100010111110001001000;
		#400 //8.808989e-38 * -960501900000.0 = -8.461051e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101011111101100111110101110000;
		b = 32'b10100110010101001001011110110111;
		correct = 32'b10010010110011001011000111110101;
		#400 //1.7514167e-12 * -7.3757887e-16 = -1.291808e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010001010010010110110100010;
		b = 32'b00111000001100111100000110100101;
		correct = 32'b10110010111011011001010111000001;
		#400 //-0.0006453638 * 4.285727e-05 = -2.7658531e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010101101011000010000101101011;
		b = 32'b11010011011101011100000101100110;
		correct = 32'b00101001101001010011111000000101;
		#400 //-6.952297e-26 * -1055511700000.0 = 7.3382306e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110001101110011111000011010100;
		b = 32'b10101000011110110101000111011101;
		correct = 32'b00011010101101101000101010010110;
		#400 //-5.4115876e-09 * -1.395105e-14 = 7.5497333e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101100010110011100100001010111;
		b = 32'b10011011010000101111111001000000;
		correct = 32'b00001000001001011110001000011101;
		#400 //-3.0948766e-12 * -1.6129456e-22 = 4.9918676e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101110000000111001011111110101;
		b = 32'b00110000110010100100111001001001;
		correct = 32'b10011111010011111111110001001010;
		#400 //-2.9920916e-11 * 1.4719684e-09 = -4.4042644e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101010111111010100100110110110;
		b = 32'b00111111110111000001000101001010;
		correct = 32'b10101011010110011011110001110100;
		#400 //-4.4992975e-13 * 1.7192776 = -7.735542e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101111000101001001001100010010;
		b = 32'b11110010010001011100011100100111;
		correct = 32'b01100001111001011001000110000100;
		#400 //-1.3512771e-10 * -3.9173957e+30 = 5.2934874e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000001001110100111000010010110;
		b = 32'b11110000000111101111010011111001;
		correct = 32'b01110001111001111000011111001010;
		#400 //-11.652487 * -1.9677914e+29 = 2.2929663e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010001110010101101110100000000;
		b = 32'b10000101001001110000010110001110;
		correct = 32'b00010111100001000101101010010010;
		#400 //-108911395000.0 * -7.8533225e-36 = 8.553163e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111111001111101001000110010100;
		b = 32'b10101111100110110000110010001010;
		correct = 32'b01101111011001101101011011110100;
		#400 //-2.533092e+38 * -2.8203245e-10 = 7.1441415e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000111100011110001110000001110;
		b = 32'b00111010001111000101101111101011;
		correct = 32'b11000010010100101001011111111001;
		#400 //-73272.11 * 0.00071853277 = -52.64841
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001001111101011110100110011101;
		b = 32'b01101010001000101001011010001100;
		correct = 32'b01110100100111000010111001110011;
		#400 //2014515.6 * 4.913923e+25 = 9.899175e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100001111000101011101100001101;
		b = 32'b10111110101011111011111010001001;
		correct = 32'b00100001000110111010011010011110;
		#400 //-1.5363868e-18 * -0.34325054 = 5.273656e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010011110101011001111001001101;
		b = 32'b01101101000101101100111111011101;
		correct = 32'b01000001011110111011000001101001;
		#400 //5.3924856e-27 * 2.9171277e+27 = 15.730569
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110111110010101100001100011011;
		b = 32'b01010111001001000001000110110001;
		correct = 32'b01001111100000011111001100000000;
		#400 //2.417113e-05 * 180395890000000.0 = 4360372000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100011001001000111100011001;
		b = 32'b00010010001100010001111011011110;
		correct = 32'b00010111000111100010001001111111;
		#400 //914.2359 * 5.58894e-28 = 5.1096094e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110111100101101001010101000010;
		b = 32'b11000101101001101111111100100011;
		correct = 32'b01111101110001000111010110111000;
		#400 //-6.108374e+33 * -5343.892 = 3.264249e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001101000101111011101100010011;
		b = 32'b00010101101100010000101001010101;
		correct = 32'b00100011010100011101110011110000;
		#400 //159101230.0 * 7.150603e-26 = 1.1376698e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001001001010001110001001001100;
		b = 32'b01001000011110001101111110100011;
		correct = 32'b10010010001001000010111011000010;
		#400 //-2.0328669e-33 * 254846.55 = -5.180691e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010111110011101011000101000111;
		b = 32'b00101011001110111100010111100001;
		correct = 32'b11000011100101111001101101000011;
		#400 //-454521600000000.0 * 6.671036e-13 = -303.21298
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001010101001011100110101010111;
		b = 32'b10111110000111110001000101011010;
		correct = 32'b11001001010011100000101110001100;
		#400 //5433003.5 * -0.15533963 = -843960.75
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111111010000001100010111001000;
		b = 32'b10110100111000001111111100010110;
		correct = 32'b01110100101010010110110100100101;
		#400 //-2.5623871e+38 * -4.190885e-07 = 1.073867e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001001000011010010101110001000;
		b = 32'b01110010010100010100010111100100;
		correct = 32'b00111011111001101100111000101001;
		#400 //1.6992726e-33 * 4.145079e+30 = 0.007043619
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010000100111011100010000000000;
		b = 32'b00001011001010111111001111101000;
		correct = 32'b10011100010100111111000001111000;
		#400 //-21174944000.0 * 3.3116897e-32 = -7.012484e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000100111011000110001111111000;
		b = 32'b01111000000010100101110101000001;
		correct = 32'b00111101011111111000100000000000;
		#400 //5.557514e-36 * 1.1225443e+34 = 0.06238556
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110010001001100100011101100011;
		b = 32'b11101100001100111111100100010101;
		correct = 32'b01011110111010011100101101100111;
		#400 //-9.678703e-09 * -8.702959e+26 = 8.423336e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100010100001101110100100011100;
		b = 32'b10100001100100100011100111001111;
		correct = 32'b00000100100110100001111011010010;
		#400 //-3.6567587e-18 * -9.908647e-19 = 3.623353e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101100010111010110001111101111;
		b = 32'b11100101000001111001000100110010;
		correct = 32'b11010001111010100111101010001000;
		#400 //3.1461463e-12 * -4.0012366e+22 = -125884760000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100001111111000001000101001000;
		b = 32'b00110110010111101001001000011100;
		correct = 32'b01011000110110110010011011011010;
		#400 //5.812281e+20 * 3.3165625e-06 = 1927679300000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110110001010010111010100110011;
		b = 32'b10111101100000010111100010110010;
		correct = 32'b10110100001010110110011111100111;
		#400 //2.5251181e-06 * -0.06321849 = -1.5963415e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011010001111001100111010001100;
		b = 32'b01001100011011101011001010010011;
		correct = 32'b01100111001100000000101110111010;
		#400 //1.3286099e+16 * 62573132.0 = 8.313528e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001101001100111011000100110010;
		b = 32'b11101010100001000100110010110111;
		correct = 32'b01111000001110011011101001101110;
		#400 //-188420900.0 * -7.997024e+25 = 1.5068065e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111110110110010011010110001001;
		b = 32'b00101100001011111111111100110100;
		correct = 32'b10101011100101010101010000100001;
		#400 //-0.42423657 * 2.5010662e-12 = -1.0610437e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010000011011111100111010110011;
		b = 32'b11101100011011000010111100110100;
		correct = 32'b10111101010111010011111011000101;
		#400 //4.7293674e-29 * -1.1421176e+27 = -0.05401494
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011101000100011001101010101011;
		b = 32'b00011011001100111111110010000011;
		correct = 32'b10111000110011001011110110001001;
		#400 //-6.557429e+17 * 1.4888124e-22 = -9.762782e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101100111000111011010010100100;
		b = 32'b00010110010100110101111111111101;
		correct = 32'b00000011101111000000001101000100;
		#400 //6.471783e-12 * 1.7074733e-25 = 1.1050397e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011100110001000010110110010001;
		b = 32'b11001100100010001011101111111111;
		correct = 32'b00101001110100011001000010001011;
		#400 //-1.2981971e-21 * -71688184.0 = 9.306539e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000111111011000110110011100111;
		b = 32'b00110110011101011011001010101101;
		correct = 32'b10111110111000101110100100111101;
		#400 //-121049.805 * 3.6611848e-06 = -0.44318572
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000000110000110101101111110001;
		b = 32'b11000011100100111010010010000100;
		correct = 32'b00000100111000010101011010101110;
		#400 //-1.7940904e-38 * -295.28528 = 5.297685e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010010100100111111011010100010;
		b = 32'b11100000101001011000111010110110;
		correct = 32'b10110011101111110110000011100101;
		#400 //9.337804e-28 * -9.543738e+19 = -8.9117556e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011111011010001110001110111;
		b = 32'b10000001111111010010111111100110;
		correct = 32'b00001110011010101000000101111111;
		#400 //-31078638.0 * -9.3006253e-38 = 2.8905077e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100110010111000110001110011101;
		b = 32'b10110001011000101101111111111011;
		correct = 32'b11011000010000110101000011000011;
		#400 //2.6018954e+23 * -3.3014647e-09 = -859006550000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100100001010000011011000110000;
		b = 32'b11001010000111001010101111110110;
		correct = 32'b11101110110011011110010000000110;
		#400 //1.241183e+22 * -2566909.5 = -3.1860045e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010001011001111101010111010110;
		b = 32'b10100100110000010001111010100010;
		correct = 32'b10110110101011101110001111110100;
		#400 //62232814000.0 * -8.37523e-17 = -5.2121413e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110011110000011010110010111001;
		b = 32'b01000000011010101111010100101101;
		correct = 32'b10110100101100011100000101011101;
		#400 //-9.018681e-08 * 3.6712143 = -3.310951e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110101111110010101100001111101;
		b = 32'b10100001100011001111110001101000;
		correct = 32'b01011000000010010101001000111101;
		#400 //-6.3216634e+32 * -9.55358e-19 = 603945200000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010011000011100111100010101111;
		b = 32'b00111101011011011001110101001101;
		correct = 32'b11010001000001000011110101000101;
		#400 //-611910100000.0 * 0.05801134 = -35497726000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100111001001001011110000111111;
		b = 32'b10000000100101001001001101000110;
		correct = 32'b00101000001111110011011100110011;
		#400 //-7.779406e+23 * -1.3644485e-38 = 1.0614599e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011011000110001111111001001011;
		b = 32'b11101000101011100101101100011110;
		correct = 32'b01000100010100000110011010010111;
		#400 //-1.2655312e-22 * -6.5869807e+24 = 833.60297
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110001010011101111101010001;
		b = 32'b00111101111010011110000110101111;
		correct = 32'b00111100100110110011001000000010;
		#400 //0.16589095 * 0.11419999 = 0.018944744
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100101000110101111011101100010;
		b = 32'b10101000001111101101011001101001;
		correct = 32'b00001101111001110000101011001010;
		#400 //-1.3441187e-16 * -1.05936115e-14 = 1.42390715e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100010010011110100111111110111;
		b = 32'b11000011000101000000000111000100;
		correct = 32'b10100101111011111011011101010010;
		#400 //2.8096064e-18 * -148.0069 = -4.1584114e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011110110100100100100000001100;
		b = 32'b00001100111001110000111110010001;
		correct = 32'b00101100001111011100101111001100;
		#400 //7.576187e+18 * 3.5600554e-31 = 2.6971645e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001101000101110111011111010011;
		b = 32'b01101010110000110011101111110101;
		correct = 32'b11111000011001110000011101111111;
		#400 //-158825780.0 * 1.1801184e+26 = -1.8743322e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111011011000011101001101001010;
		b = 32'b01110111001111001111110001101001;
		correct = 32'b11110011001001101011010111010011;
		#400 //-0.0034458213 * 3.833091e+33 = -1.3208147e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010100011100011010111101101001;
		b = 32'b01001010001010010101101101001010;
		correct = 32'b11011111000111111110001011111100;
		#400 //-4152120000000.0 * 2774738.5 = -1.1521048e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101010101111110100000110101010;
		b = 32'b00110000110010001010011010110111;
		correct = 32'b00011100000101011110011111011010;
		#400 //3.397398e-13 * 1.4599298e-09 = 4.9599626e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100001010110010011100000101100;
		b = 32'b01101011000001111001100001000000;
		correct = 32'b01001100111001100001101110011110;
		#400 //7.3596803e-19 * 1.6392397e+26 = 120642800.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001111011111010000110011001001;
		b = 32'b10011111100100011110011100001111;
		correct = 32'b10101111100100000011100010100011;
		#400 //4245473500.0 * -6.179214e-20 = -2.623369e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101110111011010000101001001111;
		b = 32'b00010101000000111011111110000111;
		correct = 32'b11000100011100111111101100111100;
		#400 //-3.6680205e+28 * 2.6606328e-26 = -975.92554
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110001101101111011101111101010;
		b = 32'b00110111011001010111100011111011;
		correct = 32'b11101001101001001011000111101101;
		#400 //-1.8196138e+30 * 1.3677632e-05 = -2.4888008e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110011000001000010100010000100;
		b = 32'b00101101100111100001110110100011;
		correct = 32'b00100001001000110100000010011100;
		#400 //3.0770494e-08 * 1.7975682e-11 = 5.531206e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111111010100010101011111100011;
		b = 32'b00000100101001000101011101111100;
		correct = 32'b00000100100001100110001111011000;
		#400 //0.8177473 * 3.8636556e-36 = 3.159494e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111101100101100111111001110110;
		b = 32'b11010101011110111110110000011000;
		correct = 32'b01010011100101000001100011001000;
		#400 //-0.07348339 * -17311965000000.0 = 1272141800000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100101110110101001100100010101;
		b = 32'b10100111001110000111111101110000;
		correct = 32'b01001101100111011000101011011001;
		#400 //-1.2903747e+23 * -2.5604214e-15 = 330390300.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101101101100110010010010110001;
		b = 32'b01011000110111111010101000001100;
		correct = 32'b01000111000111001000001111110101;
		#400 //2.0366238e-11 * 1967371500000000.0 = 40067.957
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000110010100011110001101011100;
		b = 32'b10000100111101101000000101010000;
		correct = 32'b00001011110010100001101010000000;
		#400 //-13432.84 * -5.7953077e-36 = 7.784744e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110101010101000111001001110101;
		b = 32'b01011110010011001110010010101010;
		correct = 32'b01010100001010100000100011111000;
		#400 //7.914271e-07 * 3.691028e+18 = 2921179600000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010000101000101111101101110010;
		b = 32'b10111111011011111010001001010010;
		correct = 32'b00010000100110001001000000010111;
		#400 //-6.4285146e-29 * -0.93607056 = 6.0175434e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110101111111111000100010001101;
		b = 32'b11010001011010010101011010010011;
		correct = 32'b11000111111010001110100110110011;
		#400 //1.9038722e-06 * -62636240000.0 = -119251.4
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000101100011111010101100110110;
		b = 32'b00111101110101010101111000111100;
		correct = 32'b11000011111011110111110010101101;
		#400 //-4597.4014 * 0.104183644 = -478.97403
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101111110011111000111101010001;
		b = 32'b10000111100110001110010001011110;
		correct = 32'b10110111111101111110110010000000;
		#400 //1.2847331e+29 * -2.300464e-34 = -2.9554823e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100111000010001110011100110100;
		b = 32'b01111110100011101000101111001100;
		correct = 32'b01100110000110000111011000000011;
		#400 //1.8999127e-15 * 9.473812e+37 = 1.7999416e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111010101101110011100001011101;
		b = 32'b10111011110101100110111001000101;
		correct = 32'b01110111000110010111100000001001;
		#400 //-4.7566675e+35 * -0.006543907 = 3.1127188e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000010111110111001111011000100;
		b = 32'b01000010110110100110000100001111;
		correct = 32'b10000110010101101010010010011001;
		#400 //-3.6972262e-37 * 109.18957 = -4.0369854e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100111000001000100010100111010;
		b = 32'b10100000001110111100000010100111;
		correct = 32'b10000111110000100000010000110111;
		#400 //1.8356208e-15 * -1.590326e-19 = -2.9192353e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100011010111010011010110101001;
		b = 32'b10100010001010001110100000100110;
		correct = 32'b01000110000100011111001111010000;
		#400 //-4.080597e+21 * -2.2891144e-18 = 9340.953
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011001011101001000101111111110;
		b = 32'b01000100010110101111101011101010;
		correct = 32'b10011110010100010010111011100111;
		#400 //-1.26427755e-23 * 875.92053 = -1.1074067e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101111101110011101000000111100;
		b = 32'b11001100010101111111111100101111;
		correct = 32'b10111100100111001100011100011011;
		#400 //3.3799263e-10 * -56622268.0 = -0.01913791
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010001100010110111101111010111;
		b = 32'b00110000100000100110110011001010;
		correct = 32'b01000010100011100010000001010011;
		#400 //74884770000.0 * 9.489665e-10 = 71.06313
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101011000100000010111001011101;
		b = 32'b10110111111001010110010101010000;
		correct = 32'b10100011100000010011001010001001;
		#400 //5.122342e-13 * -2.7346105e-05 = -1.400761e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000010100110111101010101011101;
		b = 32'b01101101001101100011100010101110;
		correct = 32'b11110000010111011101100001100001;
		#400 //-77.916725 * 3.5246746e+27 = -2.746311e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111010010101010001010000000100;
		b = 32'b01010011010011100011100011110000;
		correct = 32'b01001110001010111010010101111111;
		#400 //0.0008128288 * 885718500000.0 = 719937500.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000011110010010101010111011011;
		b = 32'b00011110110111100010000110000111;
		correct = 32'b00100011001011101011001011010010;
		#400 //402.67075 * 2.3519031e-20 = 9.4704256e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010010001101101000000011010110;
		b = 32'b01001100011100111000010111011011;
		correct = 32'b00011111001011011001101110111000;
		#400 //5.7587876e-28 * 63838060.0 = 3.6762982e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010010010101101101010001001100;
		b = 32'b00110001111001001100000010011100;
		correct = 32'b00000100101111111111011010110110;
		#400 //6.778817e-28 * 6.6575705e-09 = 4.5130452e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000000111001100001100000011110;
		b = 32'b01011001101110111011100101001110;
		correct = 32'b01011011001010001011101000101011;
		#400 //7.190444 * 6604945700000000.0 = 4.749249e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010011111011110100011000001110;
		b = 32'b11001001011110111101011111101100;
		correct = 32'b00011101111010110110001110000000;
		#400 //-6.040116e-27 * -1031550.75 = 6.2306863e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000011100001110010011111010;
		b = 32'b01010101110111011000110000110011;
		correct = 32'b11000110110100000111100110011001;
		#400 //-8.7636887e-10 * 30449278000000.0 = -26684.799
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001101110010010000010110010101;
		b = 32'b01001010111110011111001100101101;
		correct = 32'b11011001010001000100010101100010;
		#400 //-421573280.0 * 8190358.5 = -3452836400000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000110011011111100001110110001;
		b = 32'b11000011011100111111100110000111;
		correct = 32'b00001010011001001000000001110101;
		#400 //-4.5094675e-35 * -243.97472 = 1.1001961e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011100100001010010011000101110;
		b = 32'b10011111001110000011110100111111;
		correct = 32'b00111100001111111010011010011000;
		#400 //-2.998252e+17 * -3.9014177e-20 = 0.011697434
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011000100101011011010011111011;
		b = 32'b00010100111010000000100001000000;
		correct = 32'b10101110000001111011000011010111;
		#400 //-1316836300000000.0 * 2.3429267e-26 = -3.085251e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111110100100100001001101111010;
		b = 32'b10100110011100010111000010100111;
		correct = 32'b00100101100010011100010010011110;
		#400 //-0.28530484 * -8.3766344e-16 = 2.3898945e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011011100101100111011101000010;
		b = 32'b10011111100010101000001001100101;
		correct = 32'b10111011101000101101000111011011;
		#400 //8.470474e+16 * -5.866099e-20 = -0.0049688644
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110001111111111001000110011111;
		b = 32'b10010010101100101000000101001010;
		correct = 32'b11000101001100100011010001010011;
		#400 //2.5310311e+30 * -1.12652515e-27 = -2851.2703
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100101000100010100001001101101;
		b = 32'b10100011101010011011000100111010;
		correct = 32'b01001001010000001001001011010100;
		#400 //-4.287303e+22 * -1.8398075e-17 = 788781.25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110011011100111011000110001110;
		b = 32'b00111111010100001011011010110111;
		correct = 32'b11110011010001101010111000110010;
		#400 //-1.9307394e+31 * 0.815288 = -1.5741087e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100111010001010100111100010101;
		b = 32'b11000101100111001000001101101001;
		correct = 32'b01101101011100010100001011110010;
		#400 //-9.31765e+23 * -5008.4263 = 4.6666762e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011011100011001011110111111110;
		b = 32'b10101101011011111011000111000000;
		correct = 32'b10001001100000111100011100011001;
		#400 //2.3283837e-22 * -1.36250455e-11 = -3.1724333e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100100000111011001101001001000;
		b = 32'b10010100110111101100110101010101;
		correct = 32'b10111001100010010010101000110011;
		#400 //1.1629024e+22 * -2.249726e-26 = -0.00026162117
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111010100111010001101110001101;
		b = 32'b00010110100110111001010110011100;
		correct = 32'b01010001101111101111011011111110;
		#400 //4.078747e+35 * 2.5136017e-25 = 102523450000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000001001000010001100111101000;
		b = 32'b11010001001111101001110100001101;
		correct = 32'b00010010111011111110100000011111;
		#400 //-2.9589617e-38 * -51167416000.0 = 1.5140243e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011011000001010111011010011110;
		b = 32'b10101011111011001000011111010001;
		correct = 32'b00000111011101101010000001010000;
		#400 //-1.103983e-22 * -1.6806505e-12 = 1.8554095e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010011101011000001000000011010;
		b = 32'b01110111110101101010110001100100;
		correct = 32'b11001100000100000100100101010100;
		#400 //-4.343478e-27 * 8.708188e+33 = -37823824.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010000100011101010101011101111;
		b = 32'b11011111010111000100100101010101;
		correct = 32'b00110000011101011000011110000111;
		#400 //-5.627249e-29 * -1.5873312e+19 = 8.9323077e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001000100001001100011110101111;
		b = 32'b10101100001111010010110101000100;
		correct = 32'b00110101010001000011110111001101;
		#400 //-271933.47 * -2.6883643e-12 = 7.310562e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001011101101111010101110001010;
		b = 32'b00111011000110101011110011011001;
		correct = 32'b10000111010111100000100101011101;
		#400 //-7.074714e-32 * 0.0023611097 = -1.6704175e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011101111010011001110111100100;
		b = 32'b00110110011100010100100001101111;
		correct = 32'b00010100110111000010111110111101;
		#400 //6.183784e-21 * 3.595396e-06 = 2.2233153e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000110101111110101100101010001;
		b = 32'b01110111101000011100001111101101;
		correct = 32'b11111110111100011101001100111100;
		#400 //-24492.658 * 6.5619816e+33 = -1.6072037e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010101110001010011001101100101;
		b = 32'b11000111101111110001011000000010;
		correct = 32'b00011110000100110011001001001100;
		#400 //-7.964875e-26 * -97836.016 = 7.792516e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001110011101100011011110111011;
		b = 32'b01011111101100101000101010001100;
		correct = 32'b00101110101010111011100000000001;
		#400 //3.0348674e-30 * 2.5730498e+19 = 7.8088654e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011001001110101011011000111111;
		b = 32'b01110111001110101100000011010001;
		correct = 32'b11010001000010000011010100001011;
		#400 //-9.652779e-24 * 3.7878047e+33 = -36562840000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110010001011100010000011010110;
		b = 32'b11011011100100010101100011101101;
		correct = 32'b01001110010001011011101000101011;
		#400 //-1.0135599e-08 * -8.182329e+16 = 829328060.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001000101001101100011101101000;
		b = 32'b11001000001010010110111010101110;
		correct = 32'b10010001010111001100001101111101;
		#400 //1.0037642e-33 * -173498.72 = -1.7415179e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100101001011111001011001100000;
		b = 32'b01001101100001011110001001001110;
		correct = 32'b00110011001101111010100010110000;
		#400 //1.522978e-16 * 280775100.0 = 4.2761428e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000001110010110000110101111101;
		b = 32'b11001010011111101001010111100110;
		correct = 32'b01001100110010011110111001000111;
		#400 //-25.381586 * -4171129.5 = 105869880.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001101001111100111011110011111;
		b = 32'b11100000100110011110100010010011;
		correct = 32'b01101110011001010000010100010000;
		#400 //-199719410.0 * -8.872221e+19 = 1.7719547e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011000100100110101001011110110;
		b = 32'b10001010111111101110000001110000;
		correct = 32'b00100100000100101010110101111001;
		#400 //-1295876200000000.0 * -2.4543734e-32 = 3.180564e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000110010001010001000010001111;
		b = 32'b00110010000101111111000111110010;
		correct = 32'b00111000111010011110111000000110;
		#400 //12612.14 * 8.844369e-09 = 0.00011154641
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101100000000001011000111010000;
		b = 32'b00000110011111010000100001000010;
		correct = 32'b00110010111111100110011111000011;
		#400 //6.223288e+26 * 4.7590078e-35 = 2.9616677e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110001001011110111101000100;
		b = 32'b01010111001110111110100111101001;
		correct = 32'b01010101111100111001101011001001;
		#400 //0.16204554 * 206613310000000.0 = 33480765000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011101101100111110010001011011;
		b = 32'b10111110001111000000100100111101;
		correct = 32'b01011100100001000010001000110001;
		#400 //-1.6203232e+18 * -0.18362899 = 2.9753833e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100101011100110010101101110;
		b = 32'b00111100111110011100011010000110;
		correct = 32'b01000010001010100010011111100110;
		#400 //1395.1697 * 0.030490171 = 42.538963
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010011111111010101100011110;
		b = 32'b10100000100101100101101111010000;
		correct = 32'b00011011100101100010100111110101;
		#400 //-0.00097529765 * -2.5471745e-19 = 2.4842532e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101010000010011110011100000110;
		b = 32'b01010011010101100011111111111100;
		correct = 32'b01111101111001101101001100101101;
		#400 //4.1678454e+25 * 920196500000.0 = 3.8352366e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001001011010010110110100100001;
		b = 32'b00111110101100111101001100101111;
		correct = 32'b11001000101000111111011111011110;
		#400 //-956114.06 * 0.35122058 = -335806.94
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001101101001001110101001001110;
		b = 32'b11010111111110010101010111100110;
		correct = 32'b01100110001000001001111100111100;
		#400 //-345852350.0 * -548294650000000.0 = 1.89629e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000101110100100011000111100010;
		b = 32'b01101110000001011011010010111011;
		correct = 32'b00110100010110111001000010011110;
		#400 //1.9766629e-35 * 1.0344999e+28 = 2.0448576e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111001001010111011110111101001;
		b = 32'b00001011011101010100000110111100;
		correct = 32'b01000101001001001000100011011001;
		#400 //5.573341e+34 * 4.7234737e-32 = 2632.553
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110110110110011010100100001000;
		b = 32'b00100110101100000101111011000111;
		correct = 32'b11011110000101011111010011001011;
		#400 //-2.2073375e+33 * 1.2238143e-15 = -2.7013712e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011010010001010100101011010011;
		b = 32'b10110101011000000011101101001111;
		correct = 32'b01010000001011001100111100101110;
		#400 //-1.388321e+16 * -8.353281e-07 = 11597036000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001100111011111100010010110100;
		b = 32'b00010101011100010001110110111110;
		correct = 32'b10100010111000011101010000001001;
		#400 //-125707680.0 * 4.8693025e-26 = -6.1210873e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010011010111001101001111011100;
		b = 32'b01011111111101000010001001100111;
		correct = 32'b10110011110100101001011110011011;
		#400 //-2.7872359e-27 * 3.5183473e+19 = -9.806464e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001011001000010110000110010100;
		b = 32'b01111100111010101010010110101111;
		correct = 32'b01001000100100111110101110100011;
		#400 //3.1080882e-32 * 9.7468634e+36 = 302941.1
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001111110001010110101000101110;
		b = 32'b01101101100010011101100010001011;
		correct = 32'b00111101110101001001100110011111;
		#400 //1.9466599e-29 * 5.332654e+27 = 0.103808634
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100101011101100001111110100111;
		b = 32'b00011001100010010100110000100010;
		correct = 32'b00111111100001000000000000100010;
		#400 //7.2642877e+22 * 1.4196218e-23 = 1.031254
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001111001101110000111101010000;
		b = 32'b10010101111000111100111010001010;
		correct = 32'b10100101101000101110011001000101;
		#400 //3071234000.0 * -9.201043e-26 = -2.8258557e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011000111110011110000011011101;
		b = 32'b01011100010000110001011101000111;
		correct = 32'b01110101101111100110110100000001;
		#400 //2197953400000000.0 * 2.1965286e+17 = 4.8278675e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110010100010101100101011011010;
		b = 32'b01000111101010101000111110111001;
		correct = 32'b01111010101110001111000101000001;
		#400 //5.498133e+30 * 87327.445 = 4.801379e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011001010001111100100010011101;
		b = 32'b00111011011101010001101100001111;
		correct = 32'b11010101001111110100100000011100;
		#400 //-3514631000000000.0 * 0.0037400161 = -13144777000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101011101101011111100110111011;
		b = 32'b11100000001110000000100111010110;
		correct = 32'b11001100100000101101001001111100;
		#400 //1.2930138e-12 * -5.3045463e+19 = -68588510.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011100111100110000000110100001;
		b = 32'b11000000100110001011011101010010;
		correct = 32'b01011110000100001111011011111100;
		#400 //-5.4720168e+17 * -4.772378 = 2.6114534e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100101010111111100001110000001;
		b = 32'b11010101100101111111010110101110;
		correct = 32'b01111011100001001101001100001111;
		#400 //-6.6043384e+22 * -20885180000000.0 = 1.379328e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001000011111010101011101001010;
		b = 32'b10000001111110001100011100011010;
		correct = 32'b00001010111101100011000110011000;
		#400 //-259421.16 * -9.138651e-38 = 2.3707593e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000001001100101100111100110100;
		b = 32'b10000000000100010100100101011100;
		correct = 32'b10000000110000010010111111111101;
		#400 //11.175587 * -1.58752e-39 = -1.7741466e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011001000010010101010110000101;
		b = 32'b00001111001110011110000110111110;
		correct = 32'b00101000110001110110111111001110;
		#400 //2416006300000000.0 * 9.1646806e-30 = 2.2141926e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000001111111110101101001000;
		b = 32'b10011101000111000011101110000100;
		correct = 32'b00001101111010100011111111111100;
		#400 //-6.981975e-10 * -2.0677197e-21 = 1.4436767e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111011001100110011000101110;
		b = 32'b11010001010011010011001111111010;
		correct = 32'b01001001001110001010111010011010;
		#400 //-1.3732859e-05 * -55083770000.0 = 756457.6
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111110001010011000001110111001;
		b = 32'b10000111101010110100010111101111;
		correct = 32'b00000110011000101101001010010111;
		#400 //-0.16554154 * -2.5770324e-34 = 4.2660593e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101001111011100101110101011101;
		b = 32'b01101001001011111111001101011101;
		correct = 32'b01010011101000111101010001101100;
		#400 //1.0585519e-13 * 1.3294454e+25 = 1407287000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011011000101111001001110111101;
		b = 32'b10111010100100100101011011000111;
		correct = 32'b10010110001011010100101101000110;
		#400 //1.2538164e-22 * -0.0011164778 = -1.3998581e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011011110101011011001000101000;
		b = 32'b11011000000000100100000000011000;
		correct = 32'b00110100010110010111001111110010;
		#400 //-3.5353025e-22 * -572847200000000.0 = 2.025188e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100000110010100001000101010110;
		b = 32'b10001011101000001001101001100000;
		correct = 32'b00101100111111011000100101100000;
		#400 //-1.1648411e+20 * -6.1862036e-32 = 7.205944e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001000010100111110101111010111;
		b = 32'b01001100011100001110000000011011;
		correct = 32'b10010101010001110110011010011110;
		#400 //-6.377273e-34 * 63144044.0 = -4.026868e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010011001010011011000000100000;
		b = 32'b00001101001100001101100010000110;
		correct = 32'b10100000111010100111000100110111;
		#400 //-728804360000.0 * 5.449482e-31 = -3.971606e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010100100000000010010101100011;
		b = 32'b01110101100111001110100011110100;
		correct = 32'b01001010100111010001011011001001;
		#400 //1.2939444e-26 * 3.9781404e+32 = 5147492.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111011100001011001110000111111;
		b = 32'b01100111101011110111010110111010;
		correct = 32'b01100011101101110010011010000001;
		#400 //0.004077464 * 1.6571716e+24 = 6.7570573e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100011001000000000110101100000;
		b = 32'b00101011100001100110100110011110;
		correct = 32'b10001111001010000001001000010001;
		#400 //-8.67645e-18 * 9.550587e-13 = -8.286519e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001000111111111101000001101011;
		b = 32'b01100100100000001001000101001100;
		correct = 32'b00101110000000000111100101100110;
		#400 //1.5396253e-33 * 1.8973224e+22 = 2.9211654e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111100100101001000011000101001;
		b = 32'b11111101011001110010001011001000;
		correct = 32'b11111010100001100001100100111101;
		#400 //0.018130379 * -1.9202016e+37 = -3.4813984e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111101110101110110010111110;
		b = 32'b11110110100100000100100011101001;
		correct = 32'b11111110110100101011010011001111;
		#400 //95705.484 * -1.4632218e+33 = -1.4003835e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010010101101101001111101101110;
		b = 32'b11100010011000001000011001110010;
		correct = 32'b11110101101000000010101101101001;
		#400 //392179420000.0 * -1.0354396e+21 = -4.060781e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001011111000000001110101001000;
		b = 32'b01001101111010110011000110101011;
		correct = 32'b01011010010011011110011001011100;
		#400 //29375120.0 * 493237600.0 = 1.4488913e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100101110110000101100010100;
		b = 32'b10100101010100111000100111000000;
		correct = 32'b10101010100110101000111011000111;
		#400 //1496.3462 * -1.8348004e-16 = -2.7454967e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100111010001010100100111001000;
		b = 32'b00101010001100000111001010001011;
		correct = 32'b10010010000001111111101011111111;
		#400 //-2.7379239e-15 * 1.567168e-13 = -4.2907865e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110010101000111110110110011010;
		b = 32'b00011110011100010010100000011100;
		correct = 32'b01010001100110100110110001011101;
		#400 //6.4938623e+30 * 1.2766728e-20 = 82905375000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010011000001011011111111110111;
		b = 32'b10101101010000111101000111110000;
		correct = 32'b10000000110011001001110111010001;
		#400 //1.6881606e-27 * -1.1131082e-11 = -1.8791055e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001010001110100100011011100001;
		b = 32'b11001001101011110010101010010110;
		correct = 32'b01010100011111101110101011100001;
		#400 //-3051960.2 * -1434962.8 = 4379449200000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010101000011100001001110011100;
		b = 32'b01011110111000001010111110011100;
		correct = 32'b11110100011110010110010100111101;
		#400 //-9763430000000.0 * 8.0951654e+18 = -7.9036577e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100001000110101010110000101000;
		b = 32'b01010001010001111110011100001001;
		correct = 32'b00110010111100011000111011010100;
		#400 //5.2405076e-19 * 53660914000.0 = 2.8121043e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010111010011111010111000000001;
		b = 32'b10001011110011101110100101000011;
		correct = 32'b00100011101001111101101101000001;
		#400 //-228346250000000.0 * -7.9699287e-32 = 1.8199034e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100111110110011001101000011;
		b = 32'b11100011101010110111111101100010;
		correct = 32'b11101001001010000100100000111100;
		#400 //2009.6019 * -6.327144e+21 = -1.2715041e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100111101000010111011000010110;
		b = 32'b10110010111111110000100000100011;
		correct = 32'b01011011001000001101100111000010;
		#400 //-1.5249586e+24 * -2.9689607e-08 = 4.5275424e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100000011001110100100101110001;
		b = 32'b10110000010100110010110101101100;
		correct = 32'b01010001001111101100101010010010;
		#400 //-6.6663905e+19 * -7.68259e-10 = 51215147000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010001111110101001110101110100;
		b = 32'b00111101010100111111001101110111;
		correct = 32'b11001111110011110111111000011111;
		#400 //-134547930000.0 * 0.051745858 = -6962298400.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110100001010000001111100010100;
		b = 32'b00101011001001111001101011101001;
		correct = 32'b00011111110111000010010000000100;
		#400 //1.5657525e-07 * 5.95453e-13 = 9.323321e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110001001101010100100101011000;
		b = 32'b10101010110000001010011100110110;
		correct = 32'b10011100100010000110110101101011;
		#400 //2.6380658e-09 * -3.4222077e-13 = -9.028009e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111010011010111010000000010111;
		b = 32'b00001001100100110111010100000000;
		correct = 32'b11000100100001111011100010011101;
		#400 //-3.058592e+35 * 3.549899e-33 = -1085.7692
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110101011001111110100100011101;
		b = 32'b00011101011010110011010100100101;
		correct = 32'b01010011010101010001001100100010;
		#400 //2.9398161e+32 * 3.1129466e-21 = 915149000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010001111010011001001100101110;
		b = 32'b01001001001100111001101011100010;
		correct = 32'b01011011101000111101111100111010;
		#400 //125399580000.0 * 735662.1 = 9.225172e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001110101110000001110100111001;
		b = 32'b11011010011101001110101000011000;
		correct = 32'b00101001101100000010010000110110;
		#400 //-4.5387642e-30 * -1.7234321e+16 = 7.822252e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110000000000101110011101111001;
		b = 32'b01011111100111000001110001100110;
		correct = 32'b01010000000111111010011100100110;
		#400 //4.7622667e-10 * 2.2497956e+19 = 10714126000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101010111101100010011101011001;
		b = 32'b00001101110110101011100000001000;
		correct = 32'b10111001010100100100111001110110;
		#400 //-1.4879078e+26 * 1.3479591e-30 = -0.0002005639
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011010001101010101110111100100;
		b = 32'b11100011100011101100101100001000;
		correct = 32'b00111110010010100101001111010111;
		#400 //-3.7505767e-23 * -5.268135e+21 = 0.19758545
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001100110101010010010010001010;
		b = 32'b00111110100000111010001110001010;
		correct = 32'b11001011110110110011001110111000;
		#400 //-111748180.0 * 0.25710708 = -28731248.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011100110101001000101111100101;
		b = 32'b10111110000111101100011010110111;
		correct = 32'b01011011100000111101001101010011;
		#400 //-4.786121e+17 * -0.15505491 = 7.421115e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011001110000000100100000010110;
		b = 32'b10111010110000101010100100101000;
		correct = 32'b01010101000100100011010110101110;
		#400 //-6765307000000000.0 * -0.0014851438 = 10047453000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110010101000110010110001110110;
		b = 32'b10000111011011010001110100000101;
		correct = 32'b00111010100101110010001010101000;
		#400 //-6.463975e+30 * -1.7838426e-34 = 0.0011530714
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101011110110000101110010111000;
		b = 32'b11011011000111011111010001001101;
		correct = 32'b01000111100001010111111101010110;
		#400 //-1.5373458e-12 * -4.4460183e+16 = 68350.67
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011011011000011011101101011011;
		b = 32'b10101001011111111010110010011111;
		correct = 32'b11000101011000010111000111010110;
		#400 //6.353787e+16 * -5.67711e-14 = -3607.1147
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000100100100100000000000000100;
		b = 32'b11101111010000110000011100100000;
		correct = 32'b00110100010111100111010000100111;
		#400 //-3.432445e-36 * -6.035819e+28 = 2.0717617e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101110101001010000001011001111;
		b = 32'b00111101100000100001000110010101;
		correct = 32'b01101100101001111010110110000101;
		#400 //2.553421e+28 * 0.0635101 = 1.6216803e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100110100010001010001111000101;
		b = 32'b10110000000110100011101010110101;
		correct = 32'b11010111001001001010001110110100;
		#400 //3.2263143e+23 * -5.61083e-10 = -181023000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001001001111111110110010000101;
		b = 32'b11000101101100011011100001000100;
		correct = 32'b00001111100001010011110010101101;
		#400 //-2.3102e-33 * -5687.033 = 1.3138184e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100001111101100110000110110111;
		b = 32'b01010000110000001010101000111010;
		correct = 32'b01110011001110010110110100011110;
		#400 //5.681175e+20 * 25859052000.0 = 1.469098e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111100001000001100011010110111;
		b = 32'b10010111011111111000101001111010;
		correct = 32'b10010100001000000111110011101000;
		#400 //0.009813002 * -8.2569726e-25 = -8.102569e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010111101010001010110101000110;
		b = 32'b11101110111111101000100011001010;
		correct = 32'b11000111001001111011011000001101;
		#400 //1.0900486e-24 * -3.938728e+28 = -42934.05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010000111111101110000001101110;
		b = 32'b10111100110001110011110001110011;
		correct = 32'b00001110010001100101110010100101;
		#400 //-1.00531124e-28 * -0.024320817 = 2.4449991e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010010001000001111011100000100;
		b = 32'b11111110101001001010110010001011;
		correct = 32'b01010001010011110001010101111000;
		#400 //-5.079157e-28 * -1.0944464e+38 = 55588650000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010100011001100111110111111010;
		b = 32'b01101000111111101101101001110011;
		correct = 32'b10111101111001010111010110101101;
		#400 //-1.1636877e-26 * 9.628086e+24 = -0.112040855
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001100000100101110110100100001;
		b = 32'b11011001010111001000100110111000;
		correct = 32'b10100101111111010010010110100110;
		#400 //1.1318789e-31 * -3879745000000000.0 = -4.3914016e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011110001010111011110011011011;
		b = 32'b00110010110001001010101000011101;
		correct = 32'b01010001100000111110111010110111;
		#400 //3.0937517e+18 * 2.2894762e-08 = 70830710000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111100011110010010001000011101;
		b = 32'b10010000001011000111110101000101;
		correct = 32'b10001101001001111101110011010100;
		#400 //0.015205887 * -3.4017523e-29 = -5.172666e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001110111111001111000001010100;
		b = 32'b01010010100000011100001011011001;
		correct = 32'b01100010000000000011010110011111;
		#400 //2121804300.0 * 278659900000.0 = 5.9126176e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011100011101101000100001100;
		b = 32'b01001010101010101100011000111011;
		correct = 32'b11010110101111101000101011010001;
		#400 //-18719256.0 * 5595933.5 = -104751710000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110100100011010011101100101111;
		b = 32'b10101000000000000101011100000110;
		correct = 32'b11011101000011011001101100110100;
		#400 //8.95159e+31 * -7.1242976e-15 = -6.377379e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000011100001000011101111010001;
		b = 32'b10110011000011101001001100000010;
		correct = 32'b00110111000100110100101000111011;
		#400 //-264.46732 * -3.3195654e-08 = 8.779166e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110011101010101111000111101110;
		b = 32'b10000010001011001001011100011000;
		correct = 32'b10110110011001100111111011100001;
		#400 //2.7087322e+31 * -1.2679926e-37 = -3.4346524e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110110011111110101011100110010;
		b = 32'b10010110111011011000000010011100;
		correct = 32'b10001101111011001110010000000000;
		#400 //3.8048715e-06 * -3.837058e-25 = -1.4599512e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111000100110101000011010000000;
		b = 32'b11000100011000110000010100100110;
		correct = 32'b10111101100010010000100001011111;
		#400 //7.368345e-05 * -908.08044 = -0.0669105
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111101100011001101001000010101;
		b = 32'b00000010100001100101011100111001;
		correct = 32'b11000000100100111100101111100011;
		#400 //-2.339784e+37 * 1.9739594e-37 = -4.6186385
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100101000110100011101000010100;
		b = 32'b11001101111100010010111011001010;
		correct = 32'b01110011100100010100110011011101;
		#400 //-4.5519737e+22 * -505796930.0 = 2.3023743e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101100110101000010001100011010;
		b = 32'b11010000110010110001011010100000;
		correct = 32'b00111110001010000100101010010101;
		#400 //-6.0292995e-12 * -27258060000.0 = 0.16434701
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111010111100010011110101111010;
		b = 32'b00011100000100000001110010010100;
		correct = 32'b00010111100001111100110110000011;
		#400 //0.0018405162 * 4.768254e-22 = 8.776049e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011100010001100111000001110100;
		b = 32'b10101110011010001011110010000111;
		correct = 32'b00001011001101000110100000001100;
		#400 //-6.5658047e-22 * -5.291814e-11 = 3.4745015e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111100000010101011110101110100;
		b = 32'b00010010100101000001101011111000;
		correct = 32'b01001111001000001000100001001001;
		#400 //2.881518e+36 * 9.346761e-28 = 2693286100.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110111110110010000110101010001;
		b = 32'b10010110000100100100111001111010;
		correct = 32'b01001110011110000001100001000011;
		#400 //-8.804676e+33 * -1.1818549e-25 = 1040584900.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011100010000110100011011000011;
		b = 32'b01101011110010110110000001100011;
		correct = 32'b11001000100110110010001010100011;
		#400 //-6.4611545e-22 * 4.9173423e+26 = -317717.1
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011011111111111011000110111001;
		b = 32'b10100100110111000011111101110011;
		correct = 32'b01000001010110111111110000011011;
		#400 //-1.43943054e+17 * -9.551728e-17 = 13.749049
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010101010110111111011010111001;
		b = 32'b01011110010110001000000001101000;
		correct = 32'b11110100001110100000011010000001;
		#400 //-15115795000000.0 * 3.900146e+18 = -5.8953804e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010011001100011000101001000100;
		b = 32'b11010011000110001101100100101111;
		correct = 32'b10100110110101000000000101101110;
		#400 //2.2408711e-27 * -656478770000.0 = -1.4710843e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010001001111001011010111000001;
		b = 32'b01001100010011010110110111111111;
		correct = 32'b00011110000101110110111010100001;
		#400 //1.4886592e-28 * 53852156.0 = 8.016751e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000000110100111110010011010000;
		b = 32'b11011011010000001111100001000000;
		correct = 32'b11011100100111111011100100010111;
		#400 //6.621681 * -5.431615e+16 = -3.5966424e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000010100111100010000001110000;
		b = 32'b11110110111100010010101110011000;
		correct = 32'b00111010000101001111011101110111;
		#400 //-2.3234632e-37 * -2.4457573e+33 = 0.0005682627
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110101110000100100011111010001;
		b = 32'b11110000100011110110111000101011;
		correct = 32'b01100110110110011011001101110010;
		#400 //-1.4475028e-06 * -3.5511633e+29 = 5.1403185e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001011101011101111001101100000;
		b = 32'b11011001111111100010111001011001;
		correct = 32'b00100110001011011011010100100110;
		#400 //-6.738855e-32 * -8943200500000000.0 = 6.0266934e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010011111011101010000100001101;
		b = 32'b11111100100111100011110100111001;
		correct = 32'b11010001000100111000000001111000;
		#400 //6.0238455e-27 * -6.572997e+36 = -39594720000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011111001111010011011110100110;
		b = 32'b10000110011001000011111010001100;
		correct = 32'b10100110001010001011001111001011;
		#400 //1.3634549e+19 * -4.2927986e-35 = -5.8530374e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011111011100010001100101011110;
		b = 32'b10111011100011110010101000011100;
		correct = 32'b11011011100001101101010011010100;
		#400 //1.737302e+19 * -0.0043690335 = -7.590331e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111000101010110101110110000011;
		b = 32'b01001101011111010100010101011111;
		correct = 32'b11000110101010011000100111011010;
		#400 //-8.171333e-05 * 265573870.0 = -21700.926
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001110000101100000100111100001;
		b = 32'b00010010101000001101100110001001;
		correct = 32'b00100001001111001000101101010111;
		#400 //629307460.0 * 1.0151046e-27 = 6.388129e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100110101101100011000101110110;
		b = 32'b10100111100000111101111011111010;
		correct = 32'b00001110101110111011010000000000;
		#400 //-1.2642193e-15 * -3.6601556e-15 = 4.6272393e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010000000000110001010111101010;
		b = 32'b00011011001100110001001111011010;
		correct = 32'b10101011101101110110010011111010;
		#400 //-8797006000.0 * 1.4812947e-22 = -1.3030959e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111100101111101010011101000000;
		b = 32'b10010111011000001011001011111110;
		correct = 32'b01010100101001110101011110100101;
		#400 //-7.919429e+36 * -7.2604224e-25 = 5749840000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111100101101101000101011011010;
		b = 32'b10011110100101011001010110011001;
		correct = 32'b11011011110101010101001011111010;
		#400 //7.582514e+36 * -1.583786e-20 = -1.2009081e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000111101010111000101100011110;
		b = 32'b11010001111100011010100101001000;
		correct = 32'b00011010001000011110111101100110;
		#400 //-2.5810986e-34 * -129740900000.0 = 3.3487404e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100100100000101101010010010011;
		b = 32'b11000011000000111011011100101100;
		correct = 32'b10101000000001101010000011000111;
		#400 //5.673863e-17 * -131.71552 = -7.473357e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011101010010000010100101100111;
		b = 32'b10000100110011011111101010100111;
		correct = 32'b00100010101000010000110100100010;
		#400 //-9.014483e+17 * -4.8425456e-36 = 4.3653042e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000000111001011100100001001000;
		b = 32'b11000101100011001111001001011011;
		correct = 32'b10000110111111010000011000100001;
		#400 //2.1102176e-38 * -4510.2944 = -9.517703e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110101101100101010101111001;
		b = 32'b01110101001001001001000011011111;
		correct = 32'b11101100011010100110101111100001;
		#400 //-5.433973e-06 * 2.0861207e+32 = -1.13359234e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000110000010101001110000000010;
		b = 32'b11101101001101001000001010011111;
		correct = 32'b01110011110000110111100011010101;
		#400 //-8871.002 * -3.4915758e+27 = 3.0973775e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101100011110110110100011001100;
		b = 32'b11101000001000110011001110110000;
		correct = 32'b11010101001000000100011001111101;
		#400 //3.572742e-12 * -3.0827968e+24 = -11014038000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001010110010101100001111010111;
		b = 32'b01101000010001111101110010100111;
		correct = 32'b11110011100111100100110100000001;
		#400 //-6644203.5 * 3.775285e+24 = -2.5083762e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111101010000101000000110111111;
		b = 32'b01100000100100010001000010010000;
		correct = 32'b11011110010111000111000000100101;
		#400 //-0.047487017 * 8.3624105e+19 = -3.9710591e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010100111011111000101010000111;
		b = 32'b11001001000011110110000010101101;
		correct = 32'b00011110100001100010100011010111;
		#400 //-2.4187472e-26 * -587274.8 = 1.4204693e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111001000000010011111010010000;
		b = 32'b01101001000011100110010100101100;
		correct = 32'b11100010100011111100011110010000;
		#400 //-0.00012325705 * 1.0759077e+25 = -1.3261322e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101001011010001001000011101110;
		b = 32'b00011010001110010010101001010110;
		correct = 32'b11000100001010000011011100110010;
		#400 //-1.75722e+25 * 3.8291302e-23 = -672.8624
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100010100101110110000001100110;
		b = 32'b01011101110101110011101011111000;
		correct = 32'b11000000111111101000100110101000;
		#400 //-4.1030698e-18 * 1.9386226e+18 = -7.9543037
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110011001100011110010010010;
		b = 32'b11111100001101110111000010110111;
		correct = 32'b01110011001001001111101010101011;
		#400 //-3.4307927e-06 * -3.8099058e+36 = 1.3070997e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111000011111000111110000110101;
		b = 32'b00110110000111111010100010110011;
		correct = 32'b00101111000111010111011110000111;
		#400 //6.019716e-05 * 2.3791042e-06 = 1.4321531e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001010001111010001110100110000;
		b = 32'b11001110110101010100101100000000;
		correct = 32'b00011001100111011001000010110000;
		#400 //-9.1055085e-33 * -1789231100.0 = 1.6291858e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101100000011111001000011101011;
		b = 32'b00000000100010100100110111011000;
		correct = 32'b10101101000110110001111110001101;
		#400 //-6.94243e+26 * 1.2701224e-38 = -8.817736e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011110100111110001000000010010;
		b = 32'b01000010010000001110111100110100;
		correct = 32'b01100001011011111100000101011100;
		#400 //5.7308404e+18 * 48.233597 = 2.7641905e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110000001001110111110101010001;
		b = 32'b00010110101000001000110011011001;
		correct = 32'b00000111010100100001010011110010;
		#400 //6.093233e-10 * 2.5938282e-25 = 1.5804799e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110000100001111011100100111110;
		b = 32'b10000001100110000111001011001010;
		correct = 32'b00110010101000011010010110110001;
		#400 //-3.3603536e+29 * -5.6000696e-38 = 1.8818215e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010011010111110111001011110000;
		b = 32'b10110000110000010101010110100000;
		correct = 32'b10000100101010001100000001100100;
		#400 //2.8203226e-27 * -1.4066934e-09 = -3.9673293e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001010001110110000000100110110;
		b = 32'b11000010111011101001100000001110;
		correct = 32'b10001101101011100100101000110011;
		#400 //9.00395e-33 * -119.29698 = -1.0741441e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111101010010100111001011100;
		b = 32'b00001110010101111001001000001000;
		correct = 32'b00010110100011101001000101100011;
		#400 //86684.72 * 2.6571108e-30 = 2.303309e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110011010010110100011011000111;
		b = 32'b10011010011011010001110101010110;
		correct = 32'b11001110001111000100011111010010;
		#400 //1.6105222e+31 * -4.903415e-23 = -789705860.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011111000000111011010011011000;
		b = 32'b10100110110110101000010010000101;
		correct = 32'b11000110011000001101100001011011;
		#400 //9.490448e+18 * -1.5162708e-15 = -14390.089
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011000001011001001000011101010;
		b = 32'b01011110000010101101000001111011;
		correct = 32'b00110110101110110010010101001110;
		#400 //2.2303642e-24 * 2.5006575e+18 = 5.577377e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011010001001110000110000011111;
		b = 32'b01100001001101011000111100000110;
		correct = 32'b01111011111011001111000111001011;
		#400 //1.1754912e+16 * 2.0932291e+20 = 2.4605724e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111000101110111101111111011101;
		b = 32'b11110010010110001111001011000011;
		correct = 32'b01101011100111110011011100001011;
		#400 //-8.958553e-05 * -4.2971036e+30 = 3.8495828e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010011010011001110100010101110;
		b = 32'b11010010111111111010101110001000;
		correct = 32'b10100110110011001010010100010010;
		#400 //2.586314e-27 * -549047240000.0 = -1.4200086e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100001100010001101110010101010;
		b = 32'b01101010001001101111011100001001;
		correct = 32'b11001100001100101000011001010000;
		#400 //-9.274128e-19 * 5.046207e+25 = -46799170.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000111000010101001010111100111;
		b = 32'b01001110100010011011101010001010;
		correct = 32'b11010110000101010001111001101000;
		#400 //-35477.902 * 1155351800.0 = -40989457000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011001101101110101101000001010;
		b = 32'b10111010011011000100100000010011;
		correct = 32'b01010100101010010011101010100000;
		#400 //-6451115000000000.0 * -0.00090134254 = 5814664300000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011001101001111000000001011110;
		b = 32'b10111000100011011101001110101110;
		correct = 32'b00010010101110011001100001101001;
		#400 //-1.7319242e-23 * -6.762832e-05 = 1.1712713e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100001001011100111000001011001;
		b = 32'b00101011110101000000111001101010;
		correct = 32'b10001101100100000111111011011100;
		#400 //-5.9102184e-19 * 1.5067507e-12 = -8.905225e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001011010100110110001101110111;
		b = 32'b01001101100000001001000110101011;
		correct = 32'b00011001010101000101010000001000;
		#400 //4.071195e-32 * 269628770.0 = 1.0977113e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111011000111101010000011100011;
		b = 32'b00011110100010101100010100011110;
		correct = 32'b10011010001010111111100110111110;
		#400 //-0.0024204783 * 1.4692844e-20 = -3.556371e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011100010111101101010111110111;
		b = 32'b01010001000100000100111000111000;
		correct = 32'b10101101111110110011100011100010;
		#400 //-7.373018e-22 * 38736724000.0 = -2.8560657e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001011010110011011000110000000;
		b = 32'b10101011110000110011000111010000;
		correct = 32'b10110111101001011111110010010000;
		#400 //14266752.0 * -1.3869409e-12 = -1.9787141e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101100110111100000011011011110;
		b = 32'b11100011110010101000111101000111;
		correct = 32'b01010001001011111010110110101111;
		#400 //-6.310382e-12 * -7.473133e+21 = 47158325000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110101100111110101011110001011;
		b = 32'b10110100110011000111101101010101;
		correct = 32'b11101010111111101000110100001101;
		#400 //4.0397987e+32 * -3.8087697e-07 = -1.5386663e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111010101000110100100110111010;
		b = 32'b10000110000001011010010110010110;
		correct = 32'b10000001001010100111110111011000;
		#400 //0.0012457885 * -2.5136173e-35 = -3.1314357e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011001101011111010011110000010;
		b = 32'b10101101101101010101000010100011;
		correct = 32'b01000111111110001101000110000110;
		#400 //-6180287000000000.0 * -2.0613128e-11 = 127395.05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010110111110000010011001001101;
		b = 32'b00110010001111101011101110011011;
		correct = 32'b00001001101110001110001001000111;
		#400 //4.0090732e-25 * 1.1102112e-08 = 4.450918e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111010111111111001011111101101;
		b = 32'b00110010010010001001001110101100;
		correct = 32'b00101101110010000100001000100001;
		#400 //0.0019500233 * 1.1675109e-08 = 2.2766735e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100001101100100110000001000100;
		b = 32'b11000110100010011100101011111011;
		correct = 32'b00101000110000000000010111100110;
		#400 //-1.208723e-18 * -17637.49 = 2.131884e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010011011010111001110101001111;
		b = 32'b00110111011111111100011011111000;
		correct = 32'b01001011011010110110100011010010;
		#400 //1011956500000.0 * 1.524551e-05 = 15427794.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111000111011000101000100111;
		b = 32'b10110001001100100110011111110000;
		correct = 32'b00101000110110111001010000001011;
		#400 //-9.390095e-06 * -2.596149e-09 = 2.4378088e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011001101101010101000110011101;
		b = 32'b01100000100110010000011011101101;
		correct = 32'b11111010110110001100010101011101;
		#400 //-6379588000000000.0 * 8.821409e+19 = -5.6276956e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110000001001101011001101110111;
		b = 32'b11000010001001101001010110100000;
		correct = 32'b10110010110110001111001110011100;
		#400 //6.0645483e-10 * -41.64612 = -2.525649e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011101000011111101111100100010;
		b = 32'b10110100111011111110001110110100;
		correct = 32'b10010010100001101101000101001001;
		#400 //1.904125e-21 * -4.4682895e-07 = -8.508182e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111101000001101111100010110110;
		b = 32'b11000001111101101111000110011110;
		correct = 32'b10111111100000100011001001100010;
		#400 //0.032952033 * -30.867977 = -1.0171626
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110101001110100101000100110111;
		b = 32'b10010111110111110010110100110000;
		correct = 32'b01001101101000100110110110100010;
		#400 //-2.3618517e+32 * -1.4422444e-24 = 340636740.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111011100110011011001110001110;
		b = 32'b00110111101011100011011101100000;
		correct = 32'b10110011110100010011001010010011;
		#400 //-0.004690594 * 2.0768202e-05 = -9.74152e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101111000000100110001100011010;
		b = 32'b01010100000010111010001101110001;
		correct = 32'b01000011100011100011111000011100;
		#400 //1.1858639e-10 * 2398970200000.0 = 284.48523
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000100001110001010001011100100;
		b = 32'b10011010101000110111101100110101;
		correct = 32'b00011111011010111101000100100111;
		#400 //-738.54517 * -6.761427e-23 = 4.9936192e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101001110111011000000011001001;
		b = 32'b01010011010001110101010100011010;
		correct = 32'b01111101101011000111100010111111;
		#400 //3.3472597e+25 * 856126260000.0 = 2.865677e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111000001001110001011101110110;
		b = 32'b01101110000011000111010110110100;
		correct = 32'b01100110101101110101101101001111;
		#400 //3.9837752e-05 * 1.0867549e+28 = 4.329387e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010110101100111111010101100111;
		b = 32'b11100010001100010001011000110101;
		correct = 32'b01111001011110001111100010010001;
		#400 //-98933290000000.0 * -8.166685e+20 = 8.0795697e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100100011000100000111101011110;
		b = 32'b10010110000111001001000011011110;
		correct = 32'b10111011000010100100000101001010;
		#400 //1.6680286e+22 * -1.2647292e-25 = -0.0021096044
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110100111111011011000101000101;
		b = 32'b00000011110100000010010110000010;
		correct = 32'b10111001010011100100010100110100;
		#400 //-1.607967e+32 * 1.2233753e-36 = -0.00019671471
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000010000110100110010111011100;
		b = 32'b11110110011100110110111000000101;
		correct = 32'b10111001000100101101000100001011;
		#400 //1.1343365e-37 * -1.23433554e+33 = -0.0001400152
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101110111000011010001110011001;
		b = 32'b01011111011111001110010010111000;
		correct = 32'b01001110110111101110011010100010;
		#400 //1.0260876e-10 * 1.8222892e+19 = 1869828400.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101000011110001100100010111100;
		b = 32'b01010100010001101000010001010111;
		correct = 32'b00111101010000001110101111011101;
		#400 //1.3810293e-14 * 3410495300000.0 = 0.047099937
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110011000101101111010011001010;
		b = 32'b01000011000111000000110011010010;
		correct = 32'b11110110101110000000100101110101;
		#400 //-1.1959983e+31 * 156.05008 = -1.8663563e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111101001011101100100101100111;
		b = 32'b11010010111000100111010111010001;
		correct = 32'b11010000100110101001111000111110;
		#400 //0.04267254 * -486319620000.0 = -20752495000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111110101100100011011011000101;
		b = 32'b00000101010001111110100110001010;
		correct = 32'b11000100100010110010101100100111;
		#400 //-1.1844348e+38 * 9.3998294e-36 = -1113.3485
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001010101010001110111010111111;
		b = 32'b10101100001010110100101101000001;
		correct = 32'b00110111011000100001001001000101;
		#400 //-5535583.5 * -2.4342336e-12 = 1.3474903e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001000001111111001101000011011;
		b = 32'b11111000000100010001100111101001;
		correct = 32'b11000000110110010011001101011011;
		#400 //5.765812e-34 * -1.1772009e+34 = -6.787519
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010001111100011011011010100111;
		b = 32'b11011001000010110111111101010110;
		correct = 32'b00101011100000111011011001100111;
		#400 //-3.8135664e-28 * -2454064300000000.0 = 9.358737e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110011101011010000100011011110;
		b = 32'b00110010111110100101111001100111;
		correct = 32'b11100111001010010011101001111000;
		#400 //-2.7418433e+31 * 2.914676e-08 = -7.991585e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111001011011001110110000100001;
		b = 32'b11100110010010110100000000110110;
		correct = 32'b11100000001111000001101010101011;
		#400 //0.00022594679 * -2.3995622e+23 = -5.4217336e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101100100000001010001101011101;
		b = 32'b11001100001011101101000100010000;
		correct = 32'b00111001001011111011000000101101;
		#400 //-3.6561158e-12 * -45827136.0 = 0.00016754931
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100110010010101100011000111000;
		b = 32'b01010101101101001001001100011100;
		correct = 32'b00111100100011110000011111100101;
		#400 //7.0351465e-16 * 24817990000000.0 = 0.01745982
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010010010010101011111110100;
		b = 32'b11100110101111101011000010000101;
		correct = 32'b01100001100101011111101000011100;
		#400 //-0.00076806475 * -4.5025292e+23 = 3.458234e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001001010101100101010101101111;
		b = 32'b10111010100100101000001111110110;
		correct = 32'b11000100011101010101011001101010;
		#400 //877910.94 * -0.0011178243 = -981.3502
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010111101000101110010101100110;
		b = 32'b11111011001100010100101101101000;
		correct = 32'b01010011011000011010000100101110;
		#400 //-1.0526913e-24 * -9.20566e+35 = 969071800000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100111011110000100001011010110;
		b = 32'b00101000000110010111001010100001;
		correct = 32'b11010000000101001100111100011100;
		#400 //-1.1723798e+24 * 8.518062e-15 = -9986404000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001011011001111110100101011010;
		b = 32'b01000101101010000010000011100001;
		correct = 32'b01010001100110000100111011101100;
		#400 //15198554.0 * 5380.11 = 81769890000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011101010000011101111101100101;
		b = 32'b00011101100000010101101000110001;
		correct = 32'b00111011010000111110101110111111;
		#400 //8.731247e+17 * 3.423927e-21 = 0.0029895154
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101010001101110001110010011000;
		b = 32'b10011010100011100101101110101011;
		correct = 32'b11000101010010111010011011011100;
		#400 //5.5342114e+25 * -5.887792e-23 = -3258.4287
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001011001001000100001001101010;
		b = 32'b01000110010110100011001011111011;
		correct = 32'b00010010000011000000000101000100;
		#400 //3.1635215e-32 * 13964.745 = 4.417777e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101101110100100101010000011111;
		b = 32'b11010010010001001100101011011111;
		correct = 32'b01000000101000011010111100010101;
		#400 //-2.3911593e-11 * -211304300000.0 = 5.0526223
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111111001110110010101000010010;
		b = 32'b11110010001111011011000001101101;
		correct = 32'b11110010000010101010111100001100;
		#400 //0.7311107 * -3.757181e+30 = -2.7469152e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010100100000000001111110001100;
		b = 32'b10100000011011100110101000001000;
		correct = 32'b00110101011011101010010011001010;
		#400 //-4402280700000.0 * -2.0194467e-19 = 8.890171e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100000010101010111110000001110;
		b = 32'b10100000111000101110000010010110;
		correct = 32'b01000001101111010011001011001110;
		#400 //-6.1532743e+19 * -3.8434508e-19 = 23.649807
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100111101010011101110010001001;
		b = 32'b01110001011111011011010110011000;
		correct = 32'b01011001101010000101011101110001;
		#400 //4.7146027e-15 * 1.25630785e+30 = 5922992400000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100010100000101111010110000101;
		b = 32'b10110011011010000010100101101111;
		correct = 32'b01010110011011011000011101100101;
		#400 //-1.2078841e+21 * -5.4054393e-08 = 65291443000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011100101001010000000011110111;
		b = 32'b10100011110011110011011000000001;
		correct = 32'b11000001000001011000111010010111;
		#400 //3.7155546e+17 * -2.2465857e-17 = -8.347312
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100001100100110111010010011111;
		b = 32'b10111111111001010010010100110101;
		correct = 32'b01100010000000111111110011000001;
		#400 //-3.4000935e+20 * -1.790198 = 6.086841e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000111000111011001111010110010;
		b = 32'b11101101000110000001000111001111;
		correct = 32'b00110100101110110100001001100001;
		#400 //-1.1858004e-34 * -2.9414532e+27 = 3.487976e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011110111100110110100100011000;
		b = 32'b10100101111110110011111110010110;
		correct = 32'b10000101011011101110010010000000;
		#400 //2.5772092e-20 * -4.3584647e-16 = -1.1232675e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000101111111101001011111010001;
		b = 32'b01111010101111001100001001111101;
		correct = 32'b11000001001110111011100011101001;
		#400 //-2.3941814e-35 * 4.9004825e+35 = -11.732644
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010111011000101101001110001000;
		b = 32'b00010110000000111000001101001101;
		correct = 32'b10101101111010010000110100101010;
		#400 //-249398150000000.0 * 1.0623527e-25 = -2.649488e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010011110111101001100100010100;
		b = 32'b10010011010101001110101110001100;
		correct = 32'b10100111101110010010001110010101;
		#400 //1912101900000.0 * -2.6874295e-27 = -5.1386393e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100101011001011010011101000010;
		b = 32'b01001101110010100011101011111111;
		correct = 32'b11110011101101010110101011100111;
		#400 //-6.7781705e+22 * 424108000.0 = -2.8746764e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010100001100000001000110101010;
		b = 32'b01101110010110001110001011110011;
		correct = 32'b11000011000101010010101011111110;
		#400 //-8.889213e-27 * 1.6780782e+28 = -149.16794
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110010001110011001011111000010;
		b = 32'b10010110101110010010111101110111;
		correct = 32'b00001001100001100100000100010100;
		#400 //-1.0802923e-08 * -2.9918317e-25 = 3.2320526e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001001111100000101010011001001;
		b = 32'b00001110000111110011011101011100;
		correct = 32'b00011000100101010111100010100001;
		#400 //1968793.1 * 1.9624918e-30 = 3.86374e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110101100101110000001101000110;
		b = 32'b11000001111010100001001000110000;
		correct = 32'b10111000000010100001001110111001;
		#400 //1.1251329e-06 * -29.25888 = -3.2920132e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110110001110000011000100101100;
		b = 32'b11000010011011100101001111011110;
		correct = 32'b10111001001010110111101000001111;
		#400 //2.7446758e-06 * -59.5819 = -0.00016353301
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110110101101110101000000000010;
		b = 32'b01000001001001101100011000100010;
		correct = 32'b01111000011011101101011110000011;
		#400 //1.8590099e+33 * 10.423372 = 1.9377152e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001011011011110111011011111001;
		b = 32'b11100111011100010011000001101001;
		correct = 32'b00110011011000011001110001001001;
		#400 //-4.611923e-32 * -1.1389833e+24 = 5.2529035e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111111010111001011000111110100;
		b = 32'b11000110110100001110011111101000;
		correct = 32'b01000110101101000001100010000011;
		#400 //-0.86209035 * -26739.953 = 23052.256
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110001101110001100111011101010;
		b = 32'b10110001110111110010011010100111;
		correct = 32'b00100100001000010001100000100101;
		#400 //-5.378628e-09 * -6.4945485e-09 = 3.493176e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001010110110010001011010000110;
		b = 32'b11011101101001011010011111110010;
		correct = 32'b10101001000011000111100111101111;
		#400 //2.0904812e-32 * -1.4920969e+18 = -3.1192005e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011100010010010010100011101001;
		b = 32'b00111011100100101100011111101111;
		correct = 32'b11011000011001101010110011011111;
		#400 //-2.264858e+17 * 0.0044794003 = -1014520600000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011011111000110100101111111010;
		b = 32'b11110001011011100000000110111111;
		correct = 32'b01001101110100110101001000101111;
		#400 //-3.7603099e-22 * -1.1785527e+30 = 443172320.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010110100010000101111111110001;
		b = 32'b01011110000001010010010111010111;
		correct = 32'b00110101000011011101110000000001;
		#400 //2.2032533e-25 * 2.3985777e+18 = 5.284674e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000000000110101101001010100100;
		b = 32'b11100001101000001001101101101001;
		correct = 32'b11100010010000100100001101000111;
		#400 //2.4191065 * -3.703347e+20 = -8.9587905e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010011100010110011011000111101;
		b = 32'b11110010010011001001111100100010;
		correct = 32'b11000110010111101000101110000100;
		#400 //3.5142016e-27 * -4.0529486e+30 = -14242.879
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011010000011000011000001100011;
		b = 32'b11010011010000110110101011110110;
		correct = 32'b01101101110101100000011011011100;
		#400 //-9864925000000000.0 * -839313100000.0 = 8.2797606e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010001111101111110011111110011;
		b = 32'b11111011001101010110011010110100;
		correct = 32'b11001101101011111010101001110100;
		#400 //3.9112678e-28 * -9.418888e+35 = -368397950.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110000001110000010011101000010;
		b = 32'b00100010011001110001110110100110;
		correct = 32'b11010011001001100100000011000000;
		#400 //-2.279708e+29 * 3.1322033e-18 = -714050900000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000001100111111110110000100111;
		b = 32'b01100000001010010001010111111101;
		correct = 32'b11100010010100110100000101000100;
		#400 //-19.990309 * 4.873569e+19 = -9.742415e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011110100111111101000110101010;
		b = 32'b01110101110110110100000111011110;
		correct = 32'b01010101000010001110000101111011;
		#400 //1.6921495e-20 * 5.5588328e+32 = 9406376000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110100001011110010100101010100;
		b = 32'b01000111000110101011111110000100;
		correct = 32'b00111011110100111100001111001101;
		#400 //1.631318e-07 * 39615.516 = 0.0064625503
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000101001111100010111100100011;
		b = 32'b01110001100100011101000001001000;
		correct = 32'b10110111010110001010011011011101;
		#400 //-8.942415e-36 * 1.444068e+30 = -1.2913454e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011101110100010001101011010111;
		b = 32'b10100111111000001000011111101100;
		correct = 32'b00000110001101110110011010000010;
		#400 //-5.534959e-21 * -6.2319856e-15 = 3.4493785e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100111101000000101010011010;
		b = 32'b11011010010110110100101100100010;
		correct = 32'b11011111110100010000110010110001;
		#400 //1952.3313 * -1.5431407e+16 = -3.012722e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110111100111101110011011000011;
		b = 32'b01111010010001001011000100111011;
		correct = 32'b01110010011101000010110101011111;
		#400 //1.8942525e-05 * 2.5532121e+35 = 4.8364283e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000010101101000011101001111000;
		b = 32'b01000001010010110010111101000110;
		correct = 32'b01000100100011110000101110100101;
		#400 //90.1142 * 12.699041 = 1144.3639
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101010101000101001101000011000;
		b = 32'b00010110110111001001011100001101;
		correct = 32'b01000010000011000001110001011110;
		#400 //9.8286835e+25 * 3.5638243e-25 = 35.027702
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000011101100010010010110100010;
		b = 32'b00000110110111110110001000100111;
		correct = 32'b00001011000110101001001110110100;
		#400 //354.294 * 8.40275e-35 = 2.977044e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001010000000100000011100010101;
		b = 32'b11101110010111101101011100110000;
		correct = 32'b00111000111000100101111011100001;
		#400 //-6.260604e-33 * -1.7241454e+28 = 0.00010794192
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011110011011000010011101001100;
		b = 32'b00111101000001011000111001000100;
		correct = 32'b10011011111101100110011101001110;
		#400 //-1.2501862e-20 * 0.03260638 = -4.0764045e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101000000100000000000100101010;
		b = 32'b11110110110100110111001011101001;
		correct = 32'b01011111011011011110001100110010;
		#400 //-7.993858e-15 * -2.1443463e+33 = 1.71416e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010111100011100100110111110010;
		b = 32'b11000100110110010101010101001011;
		correct = 32'b10011100111100011001111011110111;
		#400 //9.196211e-25 * -1738.6654 = -1.5989134e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111111011110001000110000111111;
		b = 32'b00100100011001111011100111000100;
		correct = 32'b10100100011000001111101011101000;
		#400 //-0.97089 * 5.024749e-17 = -4.8784783e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101101100001010011000101101010;
		b = 32'b11001000111111000011011101101011;
		correct = 32'b01110111000000110011100101111010;
		#400 //-5.1526555e+27 * -516539.34 = 2.6615494e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011100000111101011111100001110;
		b = 32'b01101111111100100000001001000111;
		correct = 32'b11001100100101100001001000000101;
		#400 //-5.2524747e-22 * 1.4979625e+29 = -78680104.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000001010100110101110010111011;
		b = 32'b11101000011001001010110011010010;
		correct = 32'b00101010001111001100110101000110;
		#400 //-3.882111e-38 * -4.31955e+24 = 1.6768973e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011101010010111101010101001110;
		b = 32'b01111010011001101101100001101111;
		correct = 32'b11011000001101111100110111111000;
		#400 //-2.6977102e-21 * 2.9965452e+35 = -808381000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011100011110101111001011000111;
		b = 32'b00010111110100010000111101001001;
		correct = 32'b10110100110011001110111100110000;
		#400 //-2.8254272e+17 * 1.3510167e-24 = -3.8171993e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110100110010100011100011101100;
		b = 32'b11001000001001011100110001101111;
		correct = 32'b10111101100000101111100000101101;
		#400 //3.7666848e-07 * -169777.73 = -0.06394992
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011000100000001011010010100010;
		b = 32'b11100100000100011111111011010011;
		correct = 32'b10111101000100101100110011011010;
		#400 //3.3269617e-24 * -1.077256e+22 = -0.035839893
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010110111001011110001110111;
		b = 32'b01010011111111010001100101100011;
		correct = 32'b11001111010110100011110000100101;
		#400 //-0.0016840835 * 2174105300000.0 = -3661374700.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111001100011000101001101110010;
		b = 32'b10111001101011111010100101001000;
		correct = 32'b10110011110000001001001110101011;
		#400 //0.00026765052 * -0.00033504725 = -8.9675574e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011000011001101011010110010111;
		b = 32'b01101000001110111100110100000010;
		correct = 32'b11000001001010010011111101100111;
		#400 //-2.9818483e-24 * 3.547457e+24 = -10.577979
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001000100001010001111110101110;
		b = 32'b11000001110101001001110100101011;
		correct = 32'b00001010110111010001111111101110;
		#400 //-8.012094e-34 * -26.576742 = 2.1293536e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100110010101010101111111100001;
		b = 32'b01011000111010001111100101001101;
		correct = 32'b10111111110000100010111010101110;
		#400 //-7.402916e-16 * 2049259500000000.0 = -1.5170496
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010111001010110100100110101101;
		b = 32'b10111001001000100101000000100000;
		correct = 32'b11010000110110010011010001111000;
		#400 //188332920000000.0 * -0.00015479373 = -29152756000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111000000111010000000011111111;
		b = 32'b11110110100101011010110101010111;
		correct = 32'b01101111001101111001011111000111;
		#400 //-3.7432645e-05 * -1.5179062e+33 = 5.6819244e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100011111010010111010101101010;
		b = 32'b01001001111101011001000100001001;
		correct = 32'b01101110010111111111000110100010;
		#400 //8.613104e+21 * 2011681.1 = 1.7326818e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001010111111011100110010101110;
		b = 32'b01010111101110111011011001100111;
		correct = 32'b11100011001110100001100101011001;
		#400 //-8316503.0 * 412784170000000.0 = -3.432921e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011111011100000110111111100001;
		b = 32'b10111100010011110100001000101100;
		correct = 32'b00011100010000101010100010011101;
		#400 //-5.091452e-20 * -0.012650054 = 6.4407143e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001011110111110000101010000111;
		b = 32'b01000010010010111111000111111110;
		correct = 32'b00001110101100011011000000101111;
		#400 //8.5912315e-32 * 50.98632 = 4.3803527e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000101111000001001010100010010;
		b = 32'b00111100110100000001100111010111;
		correct = 32'b00000011001101101000111111001010;
		#400 //2.1119619e-35 * 0.025402946 = 5.3650055e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001000111111111011100111011110;
		b = 32'b00111010010001100110001011001101;
		correct = 32'b11000011110001100010110001110100;
		#400 //-523726.94 * 0.0007567823 = -396.3473
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001100010011011011000111110111;
		b = 32'b00111100111010011001100000111110;
		correct = 32'b10001001101110111011000101001101;
		#400 //-1.584618e-31 * 0.028514978 = -4.5185345e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100110011001110111111110000011;
		b = 32'b00011100010001001010111101010001;
		correct = 32'b10000011001100011101110000101010;
		#400 //-8.0317035e-16 * 6.507755e-22 = -5.226836e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011100110000000100111001000100;
		b = 32'b10111111010111110101110101100110;
		correct = 32'b11011100101001111100101001010110;
		#400 //4.33034e+17 * -0.8725189 = -3.7783033e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100110111101000100010111110;
		b = 32'b00110100111110010110111110111010;
		correct = 32'b00111010010110001101010000100000;
		#400 //1780.2732 * 4.6461156e-07 = 0.0008271355
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110100111001010001110100010011;
		b = 32'b00101011100100011011111100000110;
		correct = 32'b10100001000000100111000001101110;
		#400 //-4.2675728e-07 * 1.0355889e-12 = -4.4194513e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010111110010000110100010110101;
		b = 32'b11001001111111011111010001110000;
		correct = 32'b11100010010001101100111011010110;
		#400 //440704080000000.0 * -2080398.0 = -9.1683986e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000001001111111000110000010001;
		b = 32'b01101010000000111011101011111001;
		correct = 32'b11101011110001010010000100100110;
		#400 //-11.971696 * 3.981306e+25 = -4.7662985e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111100101010010101000000110000;
		b = 32'b00111010110010010101100011010001;
		correct = 32'b01111000000001010010101010110011;
		#400 //7.0329965e+36 * 0.0015361552 = 1.0803774e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111100001110100110010111001;
		b = 32'b11111011001110001011010000110110;
		correct = 32'b01110011010000110011110011000111;
		#400 //-1.612898e-05 * -9.590377e+35 = 1.5468301e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100100000000001001111101101000;
		b = 32'b00110110000010101010001001011010;
		correct = 32'b01011010100010110100111100000000;
		#400 //9.490679e+21 * 2.0658103e-06 = 1.9605942e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011111101011100111000001110101;
		b = 32'b01000010110001101001101110001000;
		correct = 32'b01100011000001110101010011110101;
		#400 //2.513935e+19 * 99.30377 = 2.4964322e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001001101100010010111100101101;
		b = 32'b01011100100101100000000000001101;
		correct = 32'b10100110110011111010001101011011;
		#400 //-4.2655564e-33 * 3.3777042e+17 = -1.4407788e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100001111001111000110001001111;
		b = 32'b00111110100001110101100001011100;
		correct = 32'b10100000111101001101010111010010;
		#400 //-1.5690308e-18 * 0.264346 = -4.1476702e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101101010000100011110001010110;
		b = 32'b11000010111101100010001011110111;
		correct = 32'b11110000101110101100000010000010;
		#400 //3.7570646e+27 * -123.06829 = -4.623755e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001000010010111110100000001101;
		b = 32'b11011000100101001110110101111111;
		correct = 32'b10100001011011010011111010100101;
		#400 //6.1360865e-34 * -1309982100000000.0 = -8.0381633e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001101000000110101001001001100;
		b = 32'b10111000001000000011110000011000;
		correct = 32'b10000101101001000110010010000110;
		#400 //4.0466553e-31 * -3.820294e-05 = -1.5459412e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000110011111110001111111000001;
		b = 32'b11001010100010100110110000100111;
		correct = 32'b00010001100010011111001011100110;
		#400 //-4.79835e-35 * -4535827.5 = 2.1764487e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000011100011011010110111001001;
		b = 32'b01101100000111001101011001010100;
		correct = 32'b10110000001011011001100100001000;
		#400 //-8.327134e-37 * 7.5841826e+26 = -6.3154504e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000011000000001100011111101010;
		b = 32'b11011111110100010100011110111000;
		correct = 32'b01100011010100101000111010010100;
		#400 //-128.78091 * -3.0160448e+19 = 3.88409e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001101000011000111101111001100;
		b = 32'b11011010100100010101101011010000;
		correct = 32'b01101000000111111000011111101000;
		#400 //-147307710.0 * -2.045686e+16 = 3.0134532e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111100001110110010010111100011;
		b = 32'b00010110100101010101000000011100;
		correct = 32'b00010011010110100100111100111011;
		#400 //0.011422607 * 2.4122804e-25 = 2.7554532e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100100000101111010101110101101;
		b = 32'b10100011110000000101001010000000;
		correct = 32'b10001000011000111110001101000101;
		#400 //3.288832e-17 * -2.0851622e-17 = -6.857748e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101100100000111010110100011111;
		b = 32'b00001000110011001000110011110101;
		correct = 32'b10110101110100100110110011101011;
		#400 //-1.2734946e+27 * 1.2310942e-33 = -1.5677919e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000001001000101101100000101010;
		b = 32'b00111010000010011101011010011110;
		correct = 32'b10111011101011110101110001100111;
		#400 //-10.177774 * 0.00052581157 = -0.0053515914
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111110000011110010010000111111;
		b = 32'b10000110001011110101000001100001;
		correct = 32'b00000100110001000000110101110001;
		#400 //-0.1397867 * -3.2972895e-35 = 4.6091723e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111001001111111000001101011110;
		b = 32'b00101111111011011111111111111011;
		correct = 32'b00101001101100100000110000011110;
		#400 //0.00018264118 * 4.3291934e-10 = 7.90689e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101001101010011110001011111111;
		b = 32'b01000000110010110111010000100110;
		correct = 32'b00101011000001110000010000010100;
		#400 //7.544485e-14 * 6.3579283 = 4.7967294e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100001110011001101100110000011;
		b = 32'b10100001100111110010000001111101;
		correct = 32'b01000011111111101010101000101111;
		#400 //-4.7235115e+20 * -1.0782859e-18 = 509.32956
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001111010101011010100010000110;
		b = 32'b01111100111110010111001100001000;
		correct = 32'b01001100110100000011000011101100;
		#400 //1.0534167e-29 * 1.036172e+37 = 109152100.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010011011010011010101000000100;
		b = 32'b10101000011111100110110011010000;
		correct = 32'b00111100011010000011101000000010;
		#400 //-1003579800000.0 * -1.4123427e-14 = 0.014173986
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110001111011101110111111010011;
		b = 32'b01000111101101010001110111111110;
		correct = 32'b01111010001010010000101110001110;
		#400 //2.3663156e+30 * 92731.984 = 2.1943313e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000110100011111110101110111110;
		b = 32'b01001100001000000110001111000001;
		correct = 32'b00010011001101000101011011010111;
		#400 //5.4137014e-35 * 42045188.0 = 2.276201e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010111000011111011000101100111;
		b = 32'b01011001000100001101011101100110;
		correct = 32'b11110000101000101001100101100010;
		#400 //-157992100000000.0 * 2548076900000000.0 = -4.02576e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111101001111001100111001111011;
		b = 32'b11000010110110100011011110111001;
		correct = 32'b11000000101000001111000011101110;
		#400 //0.046095353 * -109.10883 = -5.0294104
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000111000001111100010001001010;
		b = 32'b10011011110000011000011010110011;
		correct = 32'b00100011010011010100010011010111;
		#400 //-34756.29 * -3.201622e-22 = 1.112765e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011111011001111010001110111000;
		b = 32'b01001101100001100100001101111011;
		correct = 32'b01101101011100101111100110000011;
		#400 //1.6691387e+19 * 281571170.0 = 4.6998133e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100001010000111011010000110111;
		b = 32'b00110100010111001101001000111100;
		correct = 32'b01010110001010001100111110010111;
		#400 //2.2563131e+20 * 2.056558e-07 = 46402386000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000000101010101110000111101011;
		b = 32'b00010111010100110000100111101111;
		correct = 32'b10011000100011001101111011010110;
		#400 //-5.340078 * 6.8190315e-25 = -3.641416e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000101001100010010111101110010;
		b = 32'b10010000100101000011101100001000;
		correct = 32'b10010110010011010011000010010011;
		#400 //2834.9653 * -5.846666e-29 = -1.6575095e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111111100110101010110111110110;
		b = 32'b10001111000110011001111001001101;
		correct = 32'b10001111001110011010001100111100;
		#400 //1.2084339 * -7.57397e-30 = -9.152642e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011011010111001010100101011111;
		b = 32'b00111111100011010101000000000100;
		correct = 32'b11011011011100111001110010000011;
		#400 //-6.211072e+16 * 1.1040044 = -6.8570506e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000101001000010000011101011001;
		b = 32'b11011001000011011110000001001101;
		correct = 32'b01011110101100100111110001000110;
		#400 //-2576.4592 * -2495912000000000.0 = 6.430616e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111111011111101101010111110001;
		b = 32'b00001100011100100001001011001011;
		correct = 32'b01001100011100001111100011110011;
		#400 //3.3873476e+38 * 1.8648657e-31 = 63169484.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111001100101100011010110111010;
		b = 32'b10110011101101011101011001110001;
		correct = 32'b01101101110101010110001110011111;
		#400 //-9.749178e+34 * -8.467476e-08 = 8.2550927e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111010001010110001010001110010;
		b = 32'b00100001101110000111100111100110;
		correct = 32'b01011100011101101001000001010001;
		#400 //2.2207436e+35 * 1.2500591e-18 = 2.7760609e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101110111100011110100110001111;
		b = 32'b10010011001010110100000011010000;
		correct = 32'b11000010101000011101010001000001;
		#400 //3.7434121e+28 * -2.161519e-27 = -80.91456
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101001000000001100111001000010;
		b = 32'b00011101011001101100000110101110;
		correct = 32'b00000110111010000011010110000101;
		#400 //2.860061e-14 * 3.0540377e-21 = 8.734734e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000101110110101010110101001011;
		b = 32'b10010010010010111101110101100000;
		correct = 32'b00011000101011100010010010000100;
		#400 //-6997.6616 * -6.432837e-28 = 4.5014817e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011011011111001110001011110101;
		b = 32'b11001001110110010100100101100010;
		correct = 32'b01100101110101101010010011011111;
		#400 //-7.1181236e+16 * -1780012.2 = 1.2670347e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111000011111011101000110100100;
		b = 32'b00100101110011000100001110101111;
		correct = 32'b00011110110010101000011000101010;
		#400 //6.0515144e-05 * 3.5434223e-16 = 2.1443071e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111000001101101100001011000110;
		b = 32'b00111001110001111110001011010110;
		correct = 32'b00110010100011101011001101011001;
		#400 //4.357358e-05 * 0.00038125244 = 1.6612534e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001111110000111101000011010101;
		b = 32'b11111101000000011101101010001011;
		correct = 32'b11001101010001101010011011001011;
		#400 //1.9308924e-29 * -1.0787822e+37 = -208301230.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111100001110010010001001100000;
		b = 32'b10101101101001011001101100110110;
		correct = 32'b01101010011011111000011011001101;
		#400 //-3.8450885e+36 * -1.8827256e-11 = 7.2392462e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100111101100001110010010111100;
		b = 32'b10110110001111100100101011100000;
		correct = 32'b01011110100000110111110110000000;
		#400 //-1.6707118e+24 * -2.835579e-06 = 4.737435e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011101000000001110000011111010;
		b = 32'b00111110000000001000100101110111;
		correct = 32'b01011011100000010110101101100011;
		#400 //5.804186e+17 * 0.12552439 = 7.285669e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111001001011111111001100110111;
		b = 32'b10110000100100101111100010000011;
		correct = 32'b11101010010010100000011100000110;
		#400 //5.709906e+34 * -1.0693529e-09 = -6.1059046e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101001110001001000111011011001;
		b = 32'b00111100000111111100001011010111;
		correct = 32'b10100110011101010101010010100100;
		#400 //-8.7289286e-14 * 0.009751043 = -8.511616e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100101111101001010001011101100;
		b = 32'b11010011000111010101010010111010;
		correct = 32'b11111001100101100101100011100010;
		#400 //1.4440785e+23 * -675731340000.0 = -9.758091e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000000111010111101011011101001;
		b = 32'b10100010100011000110010011001111;
		correct = 32'b00100100000000010101011001100110;
		#400 //-7.369984 * -3.805381e-18 = 2.80456e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111001010100001000010100111111;
		b = 32'b00100011000000100110011100110100;
		correct = 32'b11011100110101000110111101110100;
		#400 //-6.766877e+34 * 7.069168e-18 = -4.783619e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011001001101010001000101101111;
		b = 32'b00010001110011000111110100000010;
		correct = 32'b00101011100100001010001001001111;
		#400 //3185383700000000.0 * 3.2262567e-28 = 1.0276865e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101110100010101110011011010111;
		b = 32'b10100101011101000010010000001100;
		correct = 32'b01010100100001000111011110010100;
		#400 //-2.1494e+28 * -2.117584e-16 = 4551535000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000001100110010101100010111000;
		b = 32'b01010010100110111101101000111001;
		correct = 32'b01010100101110101011011011011110;
		#400 //19.16832 * 334690550000.0 = 6415455400000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100110000111101010111100100101;
		b = 32'b10110000000001111100000101001110;
		correct = 32'b00010110101010000100110001011110;
		#400 //-5.5054627e-16 * -4.9387416e-10 = 2.7190058e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111111111101011110000101010100;
		b = 32'b11010010010011100100000010010100;
		correct = 32'b01111111111101011110000101010100;
		#400 //nan * -221461680000.0 = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100100011000000111001110011100;
		b = 32'b10110110101001110001010001101111;
		correct = 32'b01011011100100100111110101010101;
		#400 //-1.6561605e+22 * -4.9793666e-06 = 8.24663e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011000110111010011101111100110;
		b = 32'b01011001111110010111111100111010;
		correct = 32'b00110011010101111001110100110110;
		#400 //5.7187643e-24 * 8778394500000000.0 = 5.020157e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111101100000101110111011110000;
		b = 32'b00011000000100001100100100001000;
		correct = 32'b10010110000101000001101001110001;
		#400 //-0.0639323 * 1.8713059e-24 = -1.1963688e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010010101100010100101101011110;
		b = 32'b11111101011101011101001010000001;
		correct = 32'b01010000101010100011111011101010;
		#400 //-1.118885e-27 * -2.0422116e+37 = 22849999000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101001111001010001010101010111;
		b = 32'b00011110111010000001110100011111;
		correct = 32'b01001001010011111011010101100110;
		#400 //3.4618098e+25 * 2.4576e-20 = 850774.4
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110010101001111101011001000000;
		b = 32'b00001101100100011100110011011011;
		correct = 32'b10000000101111110010110101010001;
		#400 //-1.9538788e-08 * 8.985632e-31 = -1.7556836e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101101101010110101001100111110;
		b = 32'b01101010100000011111101011101000;
		correct = 32'b11011000101011011111100110111010;
		#400 //-1.9477416e-11 * 7.856815e+25 = -1530304600000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010000110111111000011000010100;
		b = 32'b10001110011010011000111100011111;
		correct = 32'b10011111110010111110110111111111;
		#400 //30000849000.0 * -2.8788378e-30 = -8.6367576e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111111110001000111010110100010;
		b = 32'b11011001100100101100101010010000;
		correct = 32'b01111111110001000111010110100010;
		#400 //nan * -5164758300000000.0 = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111001101011101000010111100101;
		b = 32'b01010010011111111010111100001111;
		correct = 32'b11001100101011100100111010110111;
		#400 //-0.00033287625 * 274538410000.0 = -91387320.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110110111010111110111001101;
		b = 32'b11101011100011010011010000000011;
		correct = 32'b01100010111101000101011010010100;
		#400 //-6.6009584e-06 * -3.414083e+26 = 2.2536221e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101111011101000101010110111101;
		b = 32'b01100010100011110011000100110011;
		correct = 32'b11010010100010001010101011011010;
		#400 //-2.2222131e-10 * 1.3207148e+21 = -293490980000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111100011011001000011000101001;
		b = 32'b11010010001110101110000110110111;
		correct = 32'b01001111001011001010101000000101;
		#400 //-0.014436283 * -200662700000.0 = 2896823600.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010001000101010011111110011101;
		b = 32'b01111101100010110010011010100001;
		correct = 32'b01001111001000100100000000011111;
		#400 //1.177363e-28 * 2.3120408e+37 = 2722111200.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111111100100110100100010000;
		b = 32'b10110111101000111010100000000010;
		correct = 32'b00110000000110101111011111111100;
		#400 //-2.8897572e-05 * -1.9509349e-05 = 5.637728e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110011001101001110000011111011;
		b = 32'b01011010010101001010100110111011;
		correct = 32'b11001110000101100100001000111101;
		#400 //-4.2114134e-08 * 1.4964829e+16 = -630230850.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110010101110010001110000010010;
		b = 32'b10111101000101000010101000000100;
		correct = 32'b00110000010101100100010100111000;
		#400 //-2.15496e-08 * -0.03617288 = 7.795111e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010110101110011100100101011110;
		b = 32'b11011110000101001010101010000101;
		correct = 32'b10110101010101111100100001010101;
		#400 //3.0015443e-25 * -2.6781302e+18 = -8.0385263e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111100100000100100101100010101;
		b = 32'b11100100100110000111101111111100;
		correct = 32'b11100001100110110011011101011110;
		#400 //0.015904943 * -2.2502713e+22 = -3.5790437e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000000010000010111011001000000;
		b = 32'b01001111100000011000000011110110;
		correct = 32'b10010000000001000111011001000001;
		#400 //-6.011727e-39 * 4345425000.0 = -2.612351e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011001000001110111111110011110;
		b = 32'b00111010000001010001011000101100;
		correct = 32'b10010011100011001110001000010011;
		#400 //-7.0051085e-24 * 0.0005076851 = -3.5563895e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111101001100110010111001010110;
		b = 32'b01000011101101110010011000001110;
		correct = 32'b11000001100000000011000011000010;
		#400 //-0.04374536 * 366.2973 = -16.023808
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101111101001100010110011100110;
		b = 32'b10000011000111010011110101010110;
		correct = 32'b10110011010011000010001010110011;
		#400 //1.0285758e+29 * -4.6208563e-37 = -4.752901e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000100010100010010011011000000;
		b = 32'b10101101111010110011111100011100;
		correct = 32'b00110010110000000011001000100010;
		#400 //-836.60547 * -2.6744433e-11 = 2.237454e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110011001010010000111011011111;
		b = 32'b10011011100001110000100000010011;
		correct = 32'b10001111001100100101100001011001;
		#400 //3.9361904e-08 * -2.2339094e-22 = -8.793093e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111001100000011010111110000101;
		b = 32'b01010111001111010010011010100111;
		correct = 32'b11010001001111111010010001010100;
		#400 //-0.0002473557 * 207973700000000.0 = -51443483000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101101001101011111111011100010;
		b = 32'b01011111011111101001001001011011;
		correct = 32'b01001101001101001111101011110000;
		#400 //1.0345254e-11 * 1.8343824e+19 = 189771520.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001111100110100010011010000100;
		b = 32'b11010101001000010101111110110100;
		correct = 32'b01100101010000100101011110110011;
		#400 //-5172431000.0 * -11089526000000.0 = 5.7359804e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110101011001011111111000111101;
		b = 32'b01111101111110010011001010011111;
		correct = 32'b01110011110111111110000111000100;
		#400 //8.5679113e-07 * 4.1405076e+37 = 3.5475503e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111000010100000100000001100000;
		b = 32'b01010011110101111010100011000101;
		correct = 32'b11001100101011110110111101011011;
		#400 //-4.965102e-05 * 1852498900000.0 = -91978456.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110101100000100001011010001111;
		b = 32'b10010100101011000001000100001000;
		correct = 32'b00001010101011101101111110011111;
		#400 //-9.69232e-07 * -1.737428e-26 = 1.6839707e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100001110010111010111001000000;
		b = 32'b00100110011100100000000001011110;
		correct = 32'b00001000110000001000101100000011;
		#400 //1.3801939e-18 * 8.3961114e-16 = 1.1588261e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010100001011000000100010001011;
		b = 32'b01110001101000001111010111110100;
		correct = 32'b01000110010110000101010100111110;
		#400 //8.685466e-27 * 1.5940781e+30 = 13845.311
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100000010010101111100111000011;
		b = 32'b11100000110001000011111010000010;
		correct = 32'b01000001100110111001100011001001;
		#400 //-1.7192705e-19 * -1.1312706e+20 = 19.449602
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111110111100101111110000011110;
		b = 32'b00101001001000100010100101000010;
		correct = 32'b01101000100110011110101010110100;
		#400 //1.6149112e+38 * 3.600701e-14 = 5.8148126e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000001010110101111011101011001;
		b = 32'b11000100011000110010000111101100;
		correct = 32'b01000110010000100100011001011000;
		#400 //-13.685388 * -908.53 = 12433.586
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111100000011101001110101000100;
		b = 32'b00101011110001111111110100011001;
		correct = 32'b01101000010111101101001001111110;
		#400 //2.9619835e+36 * 1.4210049e-12 = 4.208993e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110001001011011000100111011111;
		b = 32'b10000111101101011000101111000100;
		correct = 32'b10111001011101100010001001110011;
		#400 //8.593213e+29 * -2.7316e-34 = -0.00023473222
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110111110001001000000100011011;
		b = 32'b10001001001000011111111101001011;
		correct = 32'b01000001011110001011001001010000;
		#400 //-7.971162e+33 * -1.9499708e-33 = 15.543533
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010010000011000101111010000110;
		b = 32'b11011001111100110011110000011111;
		correct = 32'b01101100100001010101111010110000;
		#400 //-150720320000.0 * -8558065400000000.0 = 1.2898743e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000011101101010011010010110001;
		b = 32'b01000111000000111101100110101000;
		correct = 32'b10001011001110101010100000001110;
		#400 //-1.0650321e-36 * 33753.656 = -3.5948727e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010001100111111001011011000000;
		b = 32'b11000100001100001000011111011100;
		correct = 32'b10010110010111000001100010101011;
		#400 //2.5178684e-28 * -706.1228 = -1.7779242e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110101111000001111100010001100;
		b = 32'b00101000111100001110010111111011;
		correct = 32'b11011111010100111011001100011110;
		#400 //-5.7036896e+32 * 2.674509e-14 = -1.5254569e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011011111101111011011110111101;
		b = 32'b00110011100111111110010000011001;
		correct = 32'b11010000000110101011011111010110;
		#400 //-1.3945268e+17 * 7.445505e-08 = -10382957000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011011010101011101111001010101;
		b = 32'b01011100010011001011001111111011;
		correct = 32'b10111000001010110000001110001000;
		#400 //-1.7690786e-22 * 2.3047514e+17 = -4.0772866e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001010111101000010000111100001;
		b = 32'b00000100000111111000010101001000;
		correct = 32'b00001111100110000010000000100101;
		#400 //7999728.5 * 1.875156e-36 = 1.5000739e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000010111111010010011001111001;
		b = 32'b11101110110001101110101111000110;
		correct = 32'b10110010010001001011010011101000;
		#400 //3.719709e-37 * -3.0781532e+28 = -1.1449835e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110110000110111101100100110;
		b = 32'b00001110101001101001001011111010;
		correct = 32'b00001101111111100110010000101100;
		#400 //0.38179892 * 4.1063693e-30 = 1.5678074e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111110001100000110001111111100;
		b = 32'b00111000011010111010111010011010;
		correct = 32'b10110111001000100110010000010110;
		#400 //-0.17225641 * 5.6190976e-05 = -9.6792555e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101001100101111100011100001000;
		b = 32'b11111001101100111011010111100011;
		correct = 32'b01100011110101010001100000000010;
		#400 //-6.7402735e-14 * -1.1663878e+35 = 7.861773e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011011000011101000100100100110;
		b = 32'b01100110111010110110110101011000;
		correct = 32'b11000010100000110001010011000111;
		#400 //-1.179028e-22 * 5.5588658e+23 = -65.54058
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101111101000010011100101100101;
		b = 32'b11100100000001010011101110101001;
		correct = 32'b11010100001001111101000011001000;
		#400 //2.932651e-10 * -9.830864e+21 = -2883049200000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000011110111101010000111000010;
		b = 32'b11011000010011010110000001000101;
		correct = 32'b10011100101100101001101101000001;
		#400 //1.3085125e-36 * -903253400000000.0 = -1.1819184e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000111010110011001100010010011;
		b = 32'b00010100001001110101001101101000;
		correct = 32'b10011100000011100011100101101101;
		#400 //-55704.574 * 8.447794e-27 = -4.705808e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010101000110000011001011010101;
		b = 32'b11101000111000110111111011010101;
		correct = 32'b00111110100001110100000001111011;
		#400 //-3.0736255e-26 * -8.5945346e+24 = 0.26416382
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110100100100110000111100111;
		b = 32'b11110100100111100010000110101010;
		correct = 32'b11110011101101001101011101011001;
		#400 //0.2859032 * -1.0022775e+32 = -2.8655432e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110100010100111111111000101001;
		b = 32'b00011101001011100110011101010010;
		correct = 32'b11010010000100000110110001001111;
		#400 //-6.7183204e+31 * 2.3082124e-21 = -155073100000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100000101111100110010100001100;
		b = 32'b00010010111001100111011010000001;
		correct = 32'b10110100001010110110011011101011;
		#400 //-1.0975508e+20 * 1.4544254e-27 = -1.5963057e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011000010100100010011010010111;
		b = 32'b01111010010101101111010010111100;
		correct = 32'b01010011001100000111010100101001;
		#400 //2.7161347e-24 * 2.7902883e+35 = 757879870000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000101101111010001000100110001;
		b = 32'b11100000110100111100111101010100;
		correct = 32'b10100111000111000110111001001010;
		#400 //1.777979e-35 * -1.2210008e+20 = -2.1709137e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010011110110101010101101000101;
		b = 32'b11101010100101100100001101011001;
		correct = 32'b11111111000000000101100111100001;
		#400 //1878352600000.0 * -9.082846e+25 = -1.7060786e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100010010000010110110010001000;
		b = 32'b11011011110101100111011000111001;
		correct = 32'b10111110101000100000101000001101;
		#400 //2.6213833e-18 * -1.20731264e+17 = -0.31648293
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011110001000011000110100110001;
		b = 32'b00101100000011101010010111010011;
		correct = 32'b00001010101101000000100111101101;
		#400 //8.552467e-21 * 2.0271465e-12 = 1.7337103e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011011001111110000110000111001;
		b = 32'b00100100001000000111001000011001;
		correct = 32'b00111111111011110111100110010011;
		#400 //5.377516e+16 * 3.4791114e-17 = 1.8708977
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110011110110000101100001101100;
		b = 32'b11010101000101001101111100001011;
		correct = 32'b11001001011110111001111100111010;
		#400 //1.0074368e-07 * -10230355000000.0 = -1030643.6
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011001001100001111111111100110;
		b = 32'b11000010110011001011010010011000;
		correct = 32'b10011100100011011000100011001000;
		#400 //9.150665e-24 * -102.35272 = -9.365954e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101010101011010110101001011000;
		b = 32'b00011110110001111101111101001110;
		correct = 32'b11001010000001110110010011101111;
		#400 //-1.0482318e+26 * 2.1162301e-20 = -2218299.8
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101011100001000101011000100101;
		b = 32'b10101001001100100001011000100001;
		correct = 32'b00010101001110000001111010101100;
		#400 //-9.403074e-13 * -3.9543133e-14 = 3.71827e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001000000000010011011110100101;
		b = 32'b01010000111000010001010000001010;
		correct = 32'b00011001011000110011100000001011;
		#400 //3.8884935e-34 * 30209495000.0 = 1.1746943e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010110000010101010001001011;
		b = 32'b10010110110010010011101001011100;
		correct = 32'b00010010000101111111011101000001;
		#400 //-0.0014749853 * -3.2510131e-25 = 4.7951963e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110000011101001101001110110001;
		b = 32'b10010010010101000010100101011110;
		correct = 32'b10000011010010101110011011011110;
		#400 //8.9067514e-10 * -6.6946394e-28 = -5.9627487e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111100000100000101011000001011;
		b = 32'b00111111100101101111110100111011;
		correct = 32'b11111100001010100100001001100001;
		#400 //-2.9977436e+36 * 1.179603 = -3.5361472e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110101110101011001010110000000;
		b = 32'b10111011010010001010001100011110;
		correct = 32'b00110001101001110110010011100011;
		#400 //-1.5913247e-06 * -0.0030614804 = 4.871809e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001110000000000100110000110000;
		b = 32'b01010101100011010110001001011101;
		correct = 32'b10100100000011011011011010000100;
		#400 //-1.5813901e-30 * 19431700000000.0 = -3.0729098e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001010100010101110101011101100;
		b = 32'b01011110101101110010101111000011;
		correct = 32'b00101001110001101100101101011100;
		#400 //1.3377284e-32 * 6.599429e+18 = 8.8282436e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101010011001101001100001101011;
		b = 32'b00011001101001000001101010100110;
		correct = 32'b11000100100100111101000110100110;
		#400 //-6.969318e+25 * 1.6967966e-23 = -1182.5515
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100110100101110001001110001000;
		b = 32'b11111111111101001101001110010111;
		correct = 32'b11111111111101001101001110010111;
		#400 //-3.567188e+23 * nan = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000100001110111100010001011000;
		b = 32'b11101001110110011010101111100001;
		correct = 32'b10101110100111111010011110000000;
		#400 //2.2071901e-36 * -3.2893572e+25 = -7.260237e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001110000100101000110110110110;
		b = 32'b01001011111110101101011010011011;
		correct = 32'b11011010100011111001100100111111;
		#400 //-614690200.0 * 32877878.0 = -2.0209709e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010111010000100010010001101010;
		b = 32'b01001110001011101000000000010101;
		correct = 32'b10100110000001000101010111100010;
		#400 //-6.273074e-25 * 731907400.0 = -4.5913093e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010010100100101111001000011000;
		b = 32'b00011011010001101110100110101000;
		correct = 32'b00101110011001000101101010111011;
		#400 //315563440000.0 * 1.6453675e-22 = 5.1921783e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011110000000000101100010000000;
		b = 32'b11011000101100101111000001111001;
		correct = 32'b10110111001100110110110000110001;
		#400 //6.794565e-21 * -1573967100000000.0 = -1.0694422e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110111011011111100111000100010;
		b = 32'b10110110111101000100011111010001;
		correct = 32'b01101110111001001101001110111110;
		#400 //-4.8638274e+33 * -7.280127e-06 = 3.5409281e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010001000110111110111011001111;
		b = 32'b00000110101011011001110100111111;
		correct = 32'b00011000010100111000000001010011;
		#400 //41857905000.0 * 6.530642e-35 = 2.7335898e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100011100110011111100110001000;
		b = 32'b00001100111101100111100011101011;
		correct = 32'b00110001000101000011111010000011;
		#400 //5.680665e+21 * 3.7975076e-31 = 2.1572368e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000100101110011010100011110010;
		b = 32'b00100011001111011010100000110111;
		correct = 32'b10101000100010011000101110111001;
		#400 //-1485.2795 * 1.0281331e-17 = -1.527065e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001111000101111100110011011101;
		b = 32'b11110111111010100011111001101110;
		correct = 32'b11000111100010101110011001000111;
		#400 //7.48433e-30 * -9.50206e+33 = -71116.555
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111111001011100000100000110010;
		b = 32'b11000000110111101100011001111010;
		correct = 32'b01000000100101110111001000001001;
		#400 //-0.67981255 * -6.961728 = 4.7326703
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110101110000110101110110110100;
		b = 32'b10101010001101000000001000011010;
		correct = 32'b11100000100010010101111101111101;
		#400 //4.9531172e+32 * -1.5987941e-13 = -7.919014e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101011111000000111001100100111;
		b = 32'b00100111111101011011000100010011;
		correct = 32'b01010100010101110110100101110101;
		#400 //5.4268635e+26 * 6.8193145e-15 = 3700749000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011100011101000101100010010101;
		b = 32'b10001111110010011001011000011100;
		correct = 32'b10101100110000000110100011010100;
		#400 //2.7510917e+17 * -1.987795e-29 = -5.4686065e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110010110010101110111101001011;
		b = 32'b01001000010001110101001010101100;
		correct = 32'b10111011100111100000000110001100;
		#400 //-2.3624713e-08 * 204106.69 = -0.0048219617
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110010010010100110010010011100;
		b = 32'b00100100010110000000111110111011;
		correct = 32'b11010111001010101101000101010011;
		#400 //-4.0088065e+30 * 4.6850858e-17 = -187816020000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100001010011111000001001001101;
		b = 32'b00111011001100001000101000100010;
		correct = 32'b10011101000011110001100110001101;
		#400 //-7.030678e-19 * 0.0026937802 = -1.8939102e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111010110000000000000100100100;
		b = 32'b00100000101011011101111101111001;
		correct = 32'b11011100000000100110100001100001;
		#400 //-4.9847207e+35 * 2.9455222e-19 = -1.4682605e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000110001001101001010101111000;
		b = 32'b11101100101111101000110010110010;
		correct = 32'b01110011011101111111110011111001;
		#400 //-10661.367 * -1.8428826e+27 = 1.9647647e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110010001100000100011100011001;
		b = 32'b01100011011001010001010110111010;
		correct = 32'b11010110000111011011111010001111;
		#400 //-1.0260714e-08 * 4.22587e+21 = -43360442000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101000110001011000100001101100;
		b = 32'b00111010100001101000111100000010;
		correct = 32'b00100011110011111010011110000011;
		#400 //2.1930557e-14 * 0.0010266008 = 2.2513929e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010011110110100110001110010010;
		b = 32'b00010111011101111011001111111011;
		correct = 32'b10101011110100110100111110011100;
		#400 //-1875946800000.0 * 8.003717e-25 = -1.5014548e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110110101101101001101010011110;
		b = 32'b10000110100111010001001111101110;
		correct = 32'b00111101111000000001011000010100;
		#400 //-1.8518243e+33 * -5.908612e-35 = 0.10941711
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100000101110011110111110011110;
		b = 32'b00000000100011011000001000101100;
		correct = 32'b00100001110011011000111100001011;
		#400 //1.0718481e+20 * 1.2995502e-38 = 1.3929203e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101000111011111001001101010010;
		b = 32'b00000010110010100000110001011000;
		correct = 32'b10101100001111010001010111001100;
		#400 //-9.0509054e+24 * 2.9688317e-37 = -2.6870615e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101100111001110001101110110001;
		b = 32'b01001011011110001000101101111000;
		correct = 32'b01111000111000000110000010111100;
		#400 //2.235141e+27 * 16288632.0 = 3.640739e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101000011101001100011011011001;
		b = 32'b11000110011110111000001011111011;
		correct = 32'b00101111011100000111110000110100;
		#400 //-1.3587839e-14 * -16096.745 = 2.1871999e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101100010011010000111010101100;
		b = 32'b11101011101010010011100111100111;
		correct = 32'b01011000100001111000110100010001;
		#400 //-2.9140397e-12 * -4.091638e+26 = 1192319600000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111010011001011100100101100000;
		b = 32'b11000110101000110110100000101010;
		correct = 32'b11000001100100101010110010111000;
		#400 //0.0008765664 * -20916.082 = -18.334335
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011001100000110110100001111101;
		b = 32'b11010100010010000111011100010110;
		correct = 32'b11101110010011011100110110000101;
		#400 //4623513500000000.0 * -3443965600000.0 = -1.5923221e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000000100110001011000111001000;
		b = 32'b11101101000011100110001110111000;
		correct = 32'b01101110001010011101110000101111;
		#400 //-4.771702 * -2.754214e+27 = 1.3142288e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101111010000110111011101101110;
		b = 32'b00100000010111011011010100100010;
		correct = 32'b00010000001010010100100001100111;
		#400 //1.7777577e-10 * 1.877936e-19 = 3.338515e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110001101100110010110110111;
		b = 32'b00101110000111000101011101001000;
		correct = 32'b10100100110111101100100001010111;
		#400 //-2.717932e-06 * 3.5547815e-11 = -9.661654e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110100101011101001101000111001;
		b = 32'b11000010100111111100001000001000;
		correct = 32'b01110111110110011110110000111111;
		#400 //-1.1066744e+32 * -79.87897 = 8.8400005e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001001000001111100111010010101;
		b = 32'b10110110100010001110000110010111;
		correct = 32'b01000000000100010011101011011000;
		#400 //-556265.3 * -4.079378e-06 = 2.2692165
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001101010011001110000010001101;
		b = 32'b11101100000100001101000010011010;
		correct = 32'b01111001111001111100101010000010;
		#400 //-214829260.0 * -7.0028164e+26 = 1.5044099e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000111011011010110001011111010;
		b = 32'b01111101000010111111010110110000;
		correct = 32'b11000101000000011100100010010001;
		#400 //-1.7858985e-34 * 1.1627398e+37 = -2076.5354
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011011100100011111111101010010;
		b = 32'b10000110111010001000000000011010;
		correct = 32'b10100011000001001001100001110001;
		#400 //8.21892e+16 * -8.745693e-35 = -7.188015e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011100110011111100100010000101;
		b = 32'b01100111001000010000111101100011;
		correct = 32'b11000100100000101011100110011001;
		#400 //-1.3749944e-21 * 7.6058484e+23 = -1045.7999
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100000010010110101111100100011;
		b = 32'b10011100001001011111101010101000;
		correct = 32'b00111101000000111101101101110010;
		#400 //-5.861788e+19 * -5.4917886e-22 = 0.0321917
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100100100010001110111011000100;
		b = 32'b10111110011001110001101000000110;
		correct = 32'b11100011011101110011101010111101;
		#400 //2.0207697e+22 * -0.22568521 = -4.5605783e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000110100100001001101101010;
		b = 32'b01111000011010001010101010001100;
		correct = 32'b11101001101111101110110110001100;
		#400 //-1.5285029e-09 * 1.8876125e+34 = -2.885221e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010001001010100101011111111001;
		b = 32'b00000100100001110000111101010011;
		correct = 32'b10010110001100111011110100101101;
		#400 //-45726274000.0 * 3.175242e-36 = -1.4519198e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011101111010110101000100011110;
		b = 32'b01011100010101011111110100101100;
		correct = 32'b10111010110001001011001100110110;
		#400 //-6.2287855e-21 * 2.4093014e+17 = -0.0015007022
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100001101101101011000001111100;
		b = 32'b10111110010011101100000010011101;
		correct = 32'b11100000100100111000101101111000;
		#400 //4.2125306e+20 * -0.20190664 = -8.505379e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111111111111110010000011010011;
		b = 32'b11110101101101000101100111001011;
		correct = 32'b11110110001100111011110010010001;
		#400 //1.9931892 * -4.572435e+32 = -9.113728e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100100101010110010110101000001;
		b = 32'b01100001111010101100010001100111;
		correct = 32'b11000111000111001111101010110001;
		#400 //-7.423609e-17 * 5.413363e+20 = -40186.69
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000110101111110110001011000011;
		b = 32'b11000101101001010010110010110001;
		correct = 32'b10001100111101101111100000100010;
		#400 //7.199133e-35 * -5285.5864 = -3.805164e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010001111010000011100000001101;
		b = 32'b11100001110111111100100011101010;
		correct = 32'b01110100010010101111111100010011;
		#400 //-124671600000.0 * -5.1601266e+20 = 6.433212e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011111001110101001001001011100;
		b = 32'b10101110010000101101010101010110;
		correct = 32'b00001110000011011111111001100100;
		#400 //-3.9508098e-20 * -4.4299973e-11 = 1.7502076e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100000101001110111100010111100;
		b = 32'b00010001100110001111000111110010;
		correct = 32'b10110010110010000001101111101101;
		#400 //-9.6540815e+19 * 2.4130482e-28 = -2.3295764e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101101100011011010111110001001;
		b = 32'b10001110011111001101000101100001;
		correct = 32'b10111100100010111110110010101101;
		#400 //5.4811994e+27 * -3.116221e-30 = -0.01708063
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101001100110111100110000100100;
		b = 32'b11001111110110011010101000010010;
		correct = 32'b11111010000001000111011110001011;
		#400 //2.354344e+25 * -7303603000.0 = -1.7195195e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110100111111111001110101000;
		b = 32'b00110001110111110110011011000101;
		correct = 32'b10101001000010111001010101110110;
		#400 //-4.7669346e-06 * 6.5018377e-09 = -3.0993837e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000101010101100101001010101100;
		b = 32'b10111111001011011111100111110101;
		correct = 32'b00000101000100011010011100100010;
		#400 //-1.0077416e-35 * -0.6795953 = 6.848565e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000001100110100110011111101111;
		b = 32'b10010000101110001110000110110001;
		correct = 32'b10010010110111110000010110101000;
		#400 //19.300749 * -7.2922936e-29 = -1.4074673e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011111100011010100000000111100;
		b = 32'b01101011011101011101110011011001;
		correct = 32'b01001011100001111010100001010100;
		#400 //5.982209e-20 * 2.9722975e+26 = 17780904.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001000010101111001011111101000;
		b = 32'b11011000100101011001010101111011;
		correct = 32'b11100001011110111111001010011010;
		#400 //220767.62 * -1315754000000000.0 = -2.9047588e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010111100010011011110111011111;
		b = 32'b01111110011111111010111101110101;
		correct = 32'b11010110100010011001001010001001;
		#400 //-8.901348e-25 * 8.496604e+37 = -75631230000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110000001110110001101111110001;
		b = 32'b01001011111111000101001011010100;
		correct = 32'b11111100101110000110110000001011;
		#400 //-2.316299e+29 * 33072552.0 = -7.660592e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111010111101011010111011111101;
		b = 32'b00110010010101010110011011011111;
		correct = 32'b11101101110011001100110101010010;
		#400 //-6.3783096e+35 * 1.2421622e-08 = -7.922895e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001000001000010110111000000001;
		b = 32'b01110111101010100100000100000001;
		correct = 32'b01000000010101101011100000010100;
		#400 //4.8578484e-34 * 6.9063195e+33 = 3.3549852
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100011000100101101010110110010;
		b = 32'b00110110100110101100110000100100;
		correct = 32'b10011010001100011001001101001000;
		#400 //-7.959928e-18 * 4.6133227e-06 = -3.6721715e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111011000111010101101000111001;
		b = 32'b01100111011100011001111001000100;
		correct = 32'b11100011000101001000001100110111;
		#400 //-0.0024010076 * 1.1410098e+24 = -2.7395731e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011100011110011111000110001111;
		b = 32'b01111101101110010000100100110000;
		correct = 32'b01011010101101001010100010001001;
		#400 //8.2699396e-22 * 3.074436e+37 = 2.5425401e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000010000011001000101000010000;
		b = 32'b01111111111011001111101111001001;
		correct = 32'b01111111111011001111101111001001;
		#400 //-35.134827 * nan = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011101110111000010000010010010;
		b = 32'b10011010110000111100110100010100;
		correct = 32'b00111001001010000101110100100110;
		#400 //-1.9827298e+18 * -8.098143e-23 = 0.00016056429
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000000100101010010111111000100;
		b = 32'b01111010000100010101100101010000;
		correct = 32'b01111011001010010110100000110100;
		#400 //4.662081 * 1.8867363e+35 = 8.7961166e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110110000101011111101100010110;
		b = 32'b00100000010111010101100101000110;
		correct = 32'b11010111000000011010111000001111;
		#400 //-7.60493e+32 * 1.8748966e-19 = -142584580000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111111110011000000111000111111;
		b = 32'b10100010111011010110001011100000;
		correct = 32'b10100011001111010011100000000000;
		#400 //1.5941848 * -6.4343667e-18 = -1.0257569e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101001001000101101000000010011;
		b = 32'b01011111111010111000010001010010;
		correct = 32'b01001001100101011100100100101001;
		#400 //3.61517e-14 * 3.394156e+19 = 1227045.1
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011010110010100111001100000;
		b = 32'b01011110001000010010011101110110;
		correct = 32'b11101010000010001100101111001001;
		#400 //-14241376.0 * 2.903095e+18 = -4.1344065e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010001101110101011010111110011;
		b = 32'b01011000000110110011001101010101;
		correct = 32'b00101010011000100110001100110101;
		#400 //2.945776e-28 * 682579100000000.0 = 2.0107252e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101110111001011001011111110101;
		b = 32'b11011001001101011100001101111011;
		correct = 32'b11001000101000110000001111000001;
		#400 //1.0440707e-10 * -3197619000000000.0 = -333854.03
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111101001010110110010101010110;
		b = 32'b00100100001110010001100110001110;
		correct = 32'b11100001111101111101101010101110;
		#400 //-1.423901e+37 * 4.0137126e-17 = -5.715129e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111000001011010101001001111011;
		b = 32'b01111001001110100101100011110000;
		correct = 32'b11110001111111000101010001001000;
		#400 //-4.132323e-05 * 6.0473193e+34 = -2.4989476e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100001110110011000101101110100;
		b = 32'b11011000010110111010010000000100;
		correct = 32'b00111010101110101010010110101101;
		#400 //-1.4741405e-18 * -965989950000000.0 = 0.0014240049
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010100000011001001101111011101;
		b = 32'b00000001010011100101001111101111;
		correct = 32'b00010101111000101010011100001011;
		#400 //2415641500000.0 * 3.7896444e-38 = 9.154422e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110010001101110110110110011000;
		b = 32'b10011101010000100001101100011001;
		correct = 32'b00010000000010110001010001111000;
		#400 //-1.0676921e-08 * -2.5689695e-21 = 2.7428685e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011101100110111011001010110011;
		b = 32'b01000101100010000001011100000010;
		correct = 32'b11100011101001011000100111011011;
		#400 //-1.4024033e+18 * 4354.876 = -6.1072926e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110001011010001110110101111110;
		b = 32'b11101011110010101100000011010000;
		correct = 32'b01011101101110000111101011010101;
		#400 //-3.3895442e-09 * -4.902271e+26 = 1.6616464e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011111101011100111001001101100;
		b = 32'b01011011000101011110010011111000;
		correct = 32'b00111011010011000100100101000000;
		#400 //7.388116e-20 * 4.2191525e+16 = 0.003117159
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111100111110001110110011101010;
		b = 32'b00110000010011111111010010010111;
		correct = 32'b01101101110010100011010101100110;
		#400 //1.03399585e+37 * 7.5653744e-10 = 7.822566e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110111101110110110100010110;
		b = 32'b00001011101101100110011100010011;
		correct = 32'b10000011001100000100101100101101;
		#400 //-7.373873e-06 * 7.025894e-32 = -5.180805e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000110000010000111010110010011;
		b = 32'b01100100001000101000001000110101;
		correct = 32'b00101010101011010011111110011110;
		#400 //2.5665137e-35 * 1.199102e+22 = 3.0775117e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000001010110111110100110100101;
		b = 32'b01011010111110101001111100100011;
		correct = 32'b00011100110101110100101011011111;
		#400 //4.039158e-38 * 3.5271858e+16 = 1.424686e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101011101101010001111101000011;
		b = 32'b10011111100100011100001101100110;
		correct = 32'b00001011110011100100000111101000;
		#400 //-1.28695e-12 * -6.173315e-20 = 7.944748e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111010110001001110111110001;
		b = 32'b01111000010111111010011110100100;
		correct = 32'b11110000001111010011111101101111;
		#400 //-1.2911377e-05 * 1.8145037e+34 = -2.3427741e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111100110000001100011111110010;
		b = 32'b10100110111111001111000001011011;
		correct = 32'b11100100001111100111100111010010;
		#400 //8.007811e+36 * -1.7551161e-15 = -1.4054638e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100010110011111100101111011100;
		b = 32'b11001000001000111010101110001010;
		correct = 32'b00101011100001001101101000001010;
		#400 //-5.6323307e-18 * -167598.16 = 9.439682e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110100001001011110001001101000;
		b = 32'b01110011100101010111110110100101;
		correct = 32'b01101000010000011011110001100010;
		#400 //1.5449189e-07 * 2.3687763e+31 = 3.659567e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110111110110010010010001110111;
		b = 32'b10010010111101011110011000001101;
		correct = 32'b10001011010100001001001100001000;
		#400 //2.5885396e-05 * -1.5518386e-27 = -4.0169957e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000110000011101101010011111000;
		b = 32'b01101110100111001011001000001110;
		correct = 32'b11110101001011101101101000111110;
		#400 //-9141.242 * 2.4247458e+28 = -2.2165189e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000111100000111111000010000011;
		b = 32'b11011100001001000011110111110010;
		correct = 32'b01100100001010010100110000000010;
		#400 //-67553.02 * -1.8492002e+17 = 1.2491907e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010010111111100011101101001001;
		b = 32'b01000001110001101111100000010111;
		correct = 32'b00010101010001011001100000111011;
		#400 //1.60442685e-27 * 24.871138 = 3.9903922e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011111101110011111011101000111;
		b = 32'b11001100111110101111000010100010;
		correct = 32'b01101101001101100100101001001001;
		#400 //-2.6800515e+19 * -131564820.0 = 3.5260048e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110111101111111000111000111001;
		b = 32'b10010001011111001111101010110000;
		correct = 32'b11001001101111010100101110010101;
		#400 //7.7704165e+33 * -1.9956544e-28 = -1550706.6
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000001001101101101110110010100;
		b = 32'b11001011000101101000111100010110;
		correct = 32'b01001100110101110001100000010100;
		#400 //-11.429096 * -9867030.0 = 112771230.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100010010010010001110000011000;
		b = 32'b00101000001001000101010000101011;
		correct = 32'b10001011000000010001100000011110;
		#400 //-2.7255452e-18 * 9.12208e-15 = -2.486264e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100111011110000110011110000000;
		b = 32'b01110001001000111011011101101100;
		correct = 32'b11011001000111101101101111100001;
		#400 //-3.4473021e-15 * 8.106848e+29 = -2794675400000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101000010010111100011010000000;
		b = 32'b01011001001011000000101010010010;
		correct = 32'b01000010000010001111000111001000;
		#400 //1.13118065e-14 * 3026582400000000.0 = 34.236115
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111000000000011111011111110001;
		b = 32'b00110000110111101000100101101001;
		correct = 32'b11101001011000011111010110001100;
		#400 //-1.0544299e+34 * 1.619168e-09 = -1.7072992e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101011111010001011110101110000;
		b = 32'b01001111111011111100100011110011;
		correct = 32'b01111100010110011111111110001100;
		#400 //5.6273077e+26 * 8045848000.0 = 4.527646e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001110000110101100100110111110;
		b = 32'b01001000100011010100111011011101;
		correct = 32'b11010111001010101110000110011001;
		#400 //-649228160.0 * 289398.9 = -187885910000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010101010100110010010010111000;
		b = 32'b10110110110110010000111000001101;
		correct = 32'b10001100101100110000010110110111;
		#400 //4.2640077e-26 * -6.4687397e-06 = -2.7582756e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101101100110100111000000010111;
		b = 32'b00010111111001000110000100000111;
		correct = 32'b00000110000010011100011001011101;
		#400 //1.7557551e-11 * 1.4758648e-24 = 2.591257e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010011111000100001001100111100;
		b = 32'b11000111001000001011001111011011;
		correct = 32'b10011011100011011110101011011010;
		#400 //5.7069387e-27 * -41139.855 = -2.3478263e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101011000011000100100100011101;
		b = 32'b01110101100010011010101110111001;
		correct = 32'b11100001000101101110001001110101;
		#400 //-4.9839457e-13 * 3.4903692e+32 = -1.739581e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111001110100101011001000101011;
		b = 32'b10000111001000101111110000000011;
		correct = 32'b10000001100001100010010000101001;
		#400 //0.00040187067 * -1.2261585e-34 = -4.9275713e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001001000111100110111100101010;
		b = 32'b01101000100011011110011001001100;
		correct = 32'b10110010001011111010001110000010;
		#400 //-1.9070827e-33 * 5.360815e+24 = -1.0223518e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010110111000111100101111011000;
		b = 32'b10110111100001010111010001000110;
		correct = 32'b01001110111011011000000010111100;
		#400 //-125232320000000.0 * -1.590898e-05 = 1992318500.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100000010100110001110011011;
		b = 32'b10011100110011100111111011000100;
		correct = 32'b10100001010111110100000101011011;
		#400 //553.55634 * -1.3664705e-21 = -7.5641836e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100010000011100111011110111001;
		b = 32'b11011010011100001111011001000101;
		correct = 32'b10111101000001100001100101001011;
		#400 //1.930797e-18 * -1.6956193e+16 = -0.032738965
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010000100001011001011001111100;
		b = 32'b01000000000000100011011111010111;
		correct = 32'b00010001000001111110011100011101;
		#400 //5.269111e-29 * 2.0346582 = 1.072084e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011001101100000111011011101110;
		b = 32'b00110001010011101111100000111100;
		correct = 32'b00001011100011101010101011010000;
		#400 //1.8246009e-23 * 3.011805e-09 = 5.495342e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110010000010011110011010101010;
		b = 32'b00000011011100111011000011100001;
		correct = 32'b00110110000000110100010100111011;
		#400 //2.7314113e+30 * 7.161433e-37 = 1.9560819e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000100000110110110111110111000;
		b = 32'b11000100010100000000101111110001;
		correct = 32'b00001000111111001010010000001011;
		#400 //-1.8271461e-36 * -832.1866 = 1.5205265e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010100110100111100110111010000;
		b = 32'b11000001000101010000101111001011;
		correct = 32'b01010110011101101010000100011000;
		#400 //-7277528500000.0 * -9.315379 = 67792940000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101001011100101100111100100000;
		b = 32'b00011110100001101010011101000101;
		correct = 32'b01001000011111110110111000100011;
		#400 //1.8346136e+25 * 1.4256983e-20 = 261560.55
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110101011101000111010010101110;
		b = 32'b00111100000000111110000001110111;
		correct = 32'b11110001111110111101110000011010;
		#400 //-3.0988452e+32 * 0.008049122 = -2.4942984e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100010001011000101011010110101;
		b = 32'b11110101001011100110001101010111;
		correct = 32'b11010111111010101100101110011110;
		#400 //2.335625e-18 * -2.2106311e+32 = -516320500000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010010110110011111011111001010;
		b = 32'b01000100101000111101010110100001;
		correct = 32'b01011000000010110111111010101010;
		#400 //468082560000.0 * 1310.6759 = 613504540000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100011000011000110001011110101;
		b = 32'b10100000001110010100111101101100;
		correct = 32'b10000011110010110011111000100010;
		#400 //7.61037e-18 * -1.5696388e-19 = -1.1945533e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101011011001001000001001101000;
		b = 32'b01101010011100101011001111111010;
		correct = 32'b01010110010110001010001111101101;
		#400 //8.1182847e-13 * 7.335249e+25 = 59549640000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001110100101010011011010010001;
		b = 32'b00001011111111000001111101111111;
		correct = 32'b10011011000100101111010000010010;
		#400 //-1251690600.0 * 9.711426e-32 = -1.21557e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010010000010101011100110110010;
		b = 32'b01001110100000001001101100100110;
		correct = 32'b01100001000010110110000111011000;
		#400 //148955230000.0 * 1078825700.0 = 1.6069674e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000010101100101111100100010111;
		b = 32'b01010010111000110111011010111001;
		correct = 32'b01010110000111110000010111100000;
		#400 //89.4865 * 488474700000.0 = 43711895000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101110001001110011101010110100;
		b = 32'b01100010001111000110111001101010;
		correct = 32'b11010000111101100010111001111001;
		#400 //-3.8023543e-11 * 8.68986e+20 = -33041926000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111001101000010101000100000000;
		b = 32'b11111001000001110010101000110111;
		correct = 32'b01110011001010100101100010100010;
		#400 //-0.00030768663 * -4.386352e+34 = 1.3496218e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101111000010110011000101111001;
		b = 32'b10111111011001010101001100011010;
		correct = 32'b10101110111110010110000011100001;
		#400 //1.2659553e-10 * -0.8957993 = -1.1340418e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101111010101010111011111101000;
		b = 32'b01101010001110101111010110011110;
		correct = 32'b11011010000110111110010111101110;
		#400 //-1.9414836e-10 * 5.6505024e+25 = -1.0970358e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011101010000001000101111100010;
		b = 32'b00101101111100001000001001101101;
		correct = 32'b01001011101101001110010100111101;
		#400 //8.67152e+17 * 2.7342762e-11 = 23710330.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001001011111100010101111000001;
		b = 32'b01001100010000001110110001110101;
		correct = 32'b11010110001111111000101110010101;
		#400 //-1041084.06 * 50573780.0 = -52651555000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011011011000011001010111110111;
		b = 32'b00110001111100001101000011101000;
		correct = 32'b00001101110101000011010010101110;
		#400 //1.866002e-22 * 7.008669e-09 = 1.3078191e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010001101101001110101111100100;
		b = 32'b01111000100000010101000000001001;
		correct = 32'b11001010101101101100011011011100;
		#400 //-2.8544371e-28 * 2.0982175e+34 = -5989230.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001111100010101100101100101101;
		b = 32'b11101100111001010010100100101101;
		correct = 32'b00111100111110000111110000100100;
		#400 //-1.3686111e-29 * -2.2163077e+27 = 0.030332632
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100111110111100001011000011000;
		b = 32'b10011001100100000001001111011110;
		correct = 32'b11000001111110011111101101010011;
		#400 //2.0975458e+24 * -1.4897275e-23 = -31.247717
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101010100011011100010111010100;
		b = 32'b11000011100111101101011001110010;
		correct = 32'b01101110101011111110110110110111;
		#400 //-8.569638e+25 * -317.67535 = 2.7223628e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110010011001111001101000100011;
		b = 32'b01101000011001100010011011010010;
		correct = 32'b11011011010100000011011110011010;
		#400 //-1.3481016e-08 * 4.3474416e+24 = -5.860793e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100000010101011001010001011;
		b = 32'b11010000111101110001000010000111;
		correct = 32'b11010101100001011101101100111000;
		#400 //554.78973 * -33160444000.0 = -18397073000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101100111101000100000000110011;
		b = 32'b10000110100010010111100011011101;
		correct = 32'b00110100000000110010100110101100;
		#400 //-2.3622486e+27 * -5.1711265e-35 = 1.2215486e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100000100011101011001111110010;
		b = 32'b00101101000100010100010001011011;
		correct = 32'b00001110001000011111010000001101;
		#400 //2.4174814e-19 * 8.257474e-12 = 1.9962288e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101001011001110000010101001010;
		b = 32'b10010011110010011111110010001111;
		correct = 32'b10111101101101100100011100010001;
		#400 //1.7455428e+25 * -5.0988575e-27 = -0.089002736
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011110001101110110110100010001;
		b = 32'b10100110111111010001000111110010;
		correct = 32'b11000101101101010101001110100101;
		#400 //3.3043098e+18 * -1.7560266e-15 = -5802.4556
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111100010001001011011010101111;
		b = 32'b00110101000000011101000111001011;
		correct = 32'b01110001110001111000001010000111;
		#400 //4.0855818e+36 * 4.8361534e-07 = 1.97585e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001000101000010000110100110101;
		b = 32'b10010101001111000100001000111100;
		correct = 32'b10011110011011001101111010111100;
		#400 //329833.66 * -3.8018547e-26 = -1.2539796e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110101111001100101010010000;
		b = 32'b00111000010010101010100000110010;
		correct = 32'b10101111100101010111001111011111;
		#400 //-5.626418e-06 * 4.8317197e-05 = -2.7185273e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101111011001000111101101101010;
		b = 32'b11000001011000100010010101010000;
		correct = 32'b11110001010010011101011001000001;
		#400 //7.071178e+28 * -14.1341095 = -9.994481e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111001010000010100000000111101;
		b = 32'b01010111010000001110010000011000;
		correct = 32'b11010001000100011001110001011101;
		#400 //-0.00018429845 * 212085890000000.0 = -39087100000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010011011011100101111100001111;
		b = 32'b00111010111010010011010110011010;
		correct = 32'b00001110110110010010011001101110;
		#400 //3.008669e-27 * 0.0017792464 = 5.3531637e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001111001000010111011000000101;
		b = 32'b11011101001001111110001111010110;
		correct = 32'b10101100110100111100011101100000;
		#400 //7.9606426e-30 * -7.561093e+17 = -6.0191158e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011100000100110111111001101100;
		b = 32'b00010101101000110011011011000100;
		correct = 32'b00110010001111000001001000011001;
		#400 //1.660633e+17 * 6.592158e-26 = 1.0947155e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110100011001011011100011000000;
		b = 32'b11101111011010011101011100000001;
		correct = 32'b01100100010100011101011000010110;
		#400 //-2.1394499e-07 * -7.236993e+28 = 1.5483184e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101000011100101100010011010010;
		b = 32'b01001101110110101110110001111110;
		correct = 32'b11110110110011111001101111100000;
		#400 //-4.5857735e+24 * 459116480.0 = -2.1054042e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011010101010101110111110001110;
		b = 32'b11010000010011011100110100010101;
		correct = 32'b11101011100010010110101011000101;
		#400 //2.405707e+16 * -13811078000.0 = -3.322541e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000011111101110111011001110010;
		b = 32'b11000100010001101000011111111011;
		correct = 32'b11001000101111111110100100001110;
		#400 //494.92535 * -794.1247 = -393032.44
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100100001101001110000000101110;
		b = 32'b00101001110001101000001000010111;
		correct = 32'b11001110100011000100000101001110;
		#400 //-1.3346271e+22 * 8.8155333e-14 = -1176545000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100101001010010100110010000111;
		b = 32'b01010001100100010011100001111111;
		correct = 32'b11110111010000000001001101101010;
		#400 //-4.9968226e+22 * 77964760000.0 = -3.8957608e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001110100100101010110001010011;
		b = 32'b00000011001011100110110101111010;
		correct = 32'b10010010010001111101111110110011;
		#400 //-1230383500.0 * 5.1259677e-37 = -6.306906e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100001010010010010000100110100;
		b = 32'b10110001111100100001111101010000;
		correct = 32'b00010011101111100011100111111101;
		#400 //-6.8145393e-19 * -7.046687e-09 = 4.8019924e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010000001011111001010000101111;
		b = 32'b11011011011011110001110010111100;
		correct = 32'b01101100001000111111111100001101;
		#400 //-11782897000.0 * -6.7304113e+16 = 7.930374e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001100010111101001011001011000;
		b = 32'b00110000111101101100010011110100;
		correct = 32'b10111101110101101000111110111000;
		#400 //-58349920.0 * 1.7954833e-09 = -0.10476631
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001011000111100011000001010010;
		b = 32'b01010010101001010011011001111101;
		correct = 32'b10011110010011000010110110100001;
		#400 //-3.0466045e-32 * 354791880000.0 = -1.0809106e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110100110101010110111101100100;
		b = 32'b10011011110000111000101111111000;
		correct = 32'b11010001001000110000100010001011;
		#400 //1.3528058e+32 * -3.2350497e-22 = -43763937000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100110101110001101001110110;
		b = 32'b10100101101010011000010000010001;
		correct = 32'b10101011000011100110111101110000;
		#400 //1720.8269 * -2.9406318e-16 = -5.0603185e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010100100110101001111011111011;
		b = 32'b01001011100100010111101101001110;
		correct = 32'b11100000101011111011110100001011;
		#400 //-5312737700000.0 * 19068572.0 = -1.0130632e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010111101111000110001001011111;
		b = 32'b01010110110111100100101011101000;
		correct = 32'b01101111001000111001010001101110;
		#400 //414261370000000.0 * 122206650000000.0 = 5.0625497e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000111111010101000000110001001;
		b = 32'b11011010000010011011110011101110;
		correct = 32'b00100010011111000101100011000111;
		#400 //-3.528454e-34 * -9692451000000000.0 = 3.4199367e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101010011010000111000001110100;
		b = 32'b10011110001010100110110001001000;
		correct = 32'b11001001000110101011110011111110;
		#400 //7.025046e+25 * -9.022117e-21 = -633807.9
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001101110111110001000100000101;
		b = 32'b00010011001101101111010110010100;
		correct = 32'b00100001100111110110110000010110;
		#400 //467804320.0 * 2.3092709e-27 = 1.0802869e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110111110000101001100010000100;
		b = 32'b00101101010100111110000100100010;
		correct = 32'b01100101101000010000111011010111;
		#400 //7.893742e+33 * 1.2043951e-11 = 9.507184e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111110000100010100111011110000;
		b = 32'b10100000001100011011110001011010;
		correct = 32'b00011110110010011100010011111010;
		#400 //-0.14190269 * -1.5054803e-19 = 2.136317e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010111001010100001000011110101;
		b = 32'b01100011110100100001101001011100;
		correct = 32'b11111011100010111001001101101100;
		#400 //-186989800000000.0 * 7.7514313e+21 = -1.4494387e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100000111100000000111010111000;
		b = 32'b00100101000011000100100100010101;
		correct = 32'b10000110100000111000110010010101;
		#400 //-4.0667322e-19 * 1.2167825e-16 = -4.948329e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011001000101001101000111111001;
		b = 32'b11000110100111101011001100001111;
		correct = 32'b00100000001110001000001101011110;
		#400 //-7.693824e-24 * -20313.53 = 1.5628872e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100011010101101110100110111001;
		b = 32'b00010110111100111100101101111111;
		correct = 32'b00111010110011001010101010110001;
		#400 //3.9644447e+21 * 3.9387191e-25 = 0.0015614835
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010111000010110110110010010111;
		b = 32'b10001111111001010000111001001110;
		correct = 32'b10100111011110010111111111011011;
		#400 //153298500000000.0 * -2.2586653e-29 = -3.4625002e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111001101101110001100101111010;
		b = 32'b11011001111010101000001010011111;
		correct = 32'b01010100001001111011101010110110;
		#400 //-0.00034923461 * -8251095500000000.0 = 2881568000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100010110010011100111000111101;
		b = 32'b00000100110000010110000000011000;
		correct = 32'b00101000000110000111000000111100;
		#400 //1.8613283e+21 * 4.546233e-36 = 8.462032e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101001111101011100000100000001;
		b = 32'b00001011101100100110010011111100;
		correct = 32'b10110110001010110100000100100100;
		#400 //-3.7137283e+25 * 6.871505e-32 = -2.5518902e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110010101101011101001101011110;
		b = 32'b00011100001100011000010001110100;
		correct = 32'b01001111011111000010101001101111;
		#400 //7.202856e+30 * 5.873558e-22 = 4230639400.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000101001001100000111101100010;
		b = 32'b01110100011101110010100000000100;
		correct = 32'b11111010001000000101001011001101;
		#400 //-2656.9614 * 7.832696e+31 = -2.0811172e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000000001010101000101010000011;
		b = 32'b01001111011110000001110111000010;
		correct = 32'b11010000001001010100101000000010;
		#400 //-2.664704 * 4162699800.0 = -11092363000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111101011000000000111001110001;
		b = 32'b10110010010111010001001111111111;
		correct = 32'b00110000010000010111110111111000;
		#400 //-0.054701272 * -1.286844e-08 = 7.0392003e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101011001000110100001111000101;
		b = 32'b11110101001010001001011001001000;
		correct = 32'b01100000110101110000100010100010;
		#400 //-5.800328e-13 * -2.1370946e+32 = 1.239585e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011111100010011011000100010010;
		b = 32'b00001101100011001110110001011010;
		correct = 32'b10101101100101111001011111101011;
		#400 //-1.9843462e+19 * 8.685066e-31 = -1.7234178e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110101111101010100011010101010;
		b = 32'b00111100001001000110000010101110;
		correct = 32'b10110010100111010111110111100110;
		#400 //-1.8274488e-06 * 0.010032816 = -1.8334458e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000101110011011100110100101110;
		b = 32'b10011001001000101110101110111001;
		correct = 32'b10011111100000101111100101010111;
		#400 //6585.6475 * -8.4228075e-24 = -5.546964e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011100000000001010111110100;
		b = 32'b11001111001000110010000011111011;
		correct = 32'b01011011001000110011110011110101;
		#400 //-16788456.0 * -2736847600.0 = 4.5947444e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111001101111011100010101000110;
		b = 32'b00101010001100011110001000111010;
		correct = 32'b11100100100000111101110100011001;
		#400 //-1.2316816e+35 * 1.5799246e-13 = -1.9459642e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000000000011010000100111110111;
		b = 32'b10011101101110111101101000100111;
		correct = 32'b00011110010011101111110011101111;
		#400 //-2.2037332 * -4.9724052e-21 = 1.0957855e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111101000011011000011110100101;
		b = 32'b11100001010001101010011011110010;
		correct = 32'b11011110110110111010011001101011;
		#400 //0.03455319 * -2.2903031e+20 = -7.913728e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110111100100111010100101000011;
		b = 32'b10111101000101011001001101001111;
		correct = 32'b01110101001011001000110011111000;
		#400 //-5.989849e+33 * -0.036517438 = 2.1873395e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110100011101100010000110001101;
		b = 32'b11000010010101010001111011110101;
		correct = 32'b11110111010011001110011110101110;
		#400 //7.8002046e+31 * -53.28023 = -4.155967e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100011011001100011000110100101;
		b = 32'b11000101011011011111110011110001;
		correct = 32'b11101001010101011111111101100111;
		#400 //4.2463284e+21 * -3807.8088 = -1.6169206e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001101000101011001011100101011;
		b = 32'b11101001011111110111110101110011;
		correct = 32'b10110111000101010100101011100010;
		#400 //4.609613e-31 * -1.9304281e+25 = -8.898527e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100100000001100011101101110100;
		b = 32'b01111001101111001000110011111111;
		correct = 32'b01011110010001011011101100101111;
		#400 //2.9106977e-17 * 1.2237644e+35 = 3.5620084e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011100011101011010100100110011;
		b = 32'b00010010010100110000101000000001;
		correct = 32'b00101111010010101000010000001111;
		#400 //2.7658962e+17 * 6.659219e-28 = 1.841871e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111110011100011100110010001010;
		b = 32'b10111100001111010010110100100011;
		correct = 32'b11111011001100101010111010100100;
		#400 //8.0351494e+37 * -0.011546406 = -9.27771e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010000111010100000000100010101;
		b = 32'b11010001011010110101101100111110;
		correct = 32'b01100010110101110010001001100101;
		#400 //-31407516000.0 * -63178007000.0 = 1.9842642e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110001111110011000011101011001;
		b = 32'b11000110110101011110111110011110;
		correct = 32'b11111001010100001000011100101100;
		#400 //2.4712126e+30 * -27383.809 = -6.767121e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010000100110001011001110110001;
		b = 32'b10111001111010010111010011011001;
		correct = 32'b11001011000010110100000100111111;
		#400 //20495305000.0 * -0.0004452828 = -9126207.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110000101000010000010111011001;
		b = 32'b00010110110011000100100001101111;
		correct = 32'b11001000000000000111111000111000;
		#400 //-3.9867325e+29 * 3.300369e-25 = -131576.88
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100011111111100011011111001;
		b = 32'b11101011011010011101000011110001;
		correct = 32'b11110000011010011001110011011011;
		#400 //1023.10895 * -2.8266641e+26 = -2.8919854e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000111101011100011111101000001;
		b = 32'b00110011000010001111000111010111;
		correct = 32'b10111011001110100110110001101101;
		#400 //-89214.51 * 3.188492e-08 = -0.0028445974
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010001101011010100100010111001;
		b = 32'b01101101000001110010000111111010;
		correct = 32'b00111111001101101111000010110010;
		#400 //2.7339406e-28 * 2.613847e+27 = 0.7146102
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100101011110110011010110011000;
		b = 32'b01111110000111111010001010001010;
		correct = 32'b11100100000111001010010111001001;
		#400 //-2.1788938e-16 * 5.30478e+37 = -1.1558553e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101011011001001001010110101010;
		b = 32'b10000010100100100110110000111111;
		correct = 32'b10101110100000101011111000000010;
		#400 //2.7634186e+26 * -2.1514902e-37 = -5.945468e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101100111001111000110101110011;
		b = 32'b10100100000101100010110101101000;
		correct = 32'b10010001100001111101010111110011;
		#400 //6.581119e-12 * -3.2564526e-17 = -2.14311e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110001101101011010011010000000;
		b = 32'b10110011101010011011100000111001;
		correct = 32'b11100101111100001101101101000101;
		#400 //1.7989783e+30 * -7.903186e-08 = -1.421766e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011011011100010011000110100001;
		b = 32'b10010100110101100110010010101010;
		correct = 32'b10110000110010011111111001010100;
		#400 //6.7890037e+16 * -2.1648183e-26 = -1.4696959e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111100001001011011111001111011;
		b = 32'b10110011111011011010011011110111;
		correct = 32'b00110000100110011101110101110001;
		#400 //-0.010116215 * -1.1066543e-07 = 1.1195153e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100110110000010100111101010111;
		b = 32'b00101001111111011000000010111101;
		correct = 32'b11010001001111110110110010011111;
		#400 //-4.5644015e+23 * 1.12577895e-13 = -51385070000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111101011110010111001110010000;
		b = 32'b10000000010100010000011101111100;
		correct = 32'b00111110000111011110100110110111;
		#400 //-2.0723613e+37 * -7.44136e-39 = 0.15421186
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001111100110011001001101000011;
		b = 32'b11010101100100010100001110101111;
		correct = 32'b00100101101011100100101000000111;
		#400 //-1.5143688e-29 * -19964986000000.0 = 3.0234351e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101111000101010011000110110010;
		b = 32'b00001110010010110111001000101111;
		correct = 32'b10111101111011010010000111100111;
		#400 //-4.6173344e+28 * 2.507666e-30 = -0.11578732
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001100010011100010110100001111;
		b = 32'b01010000011101010011100011111010;
		correct = 32'b11011101010001010111111100000011;
		#400 //-54047804.0 * 16456608000.0 = -8.8944354e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111111110100000011001011110011;
		b = 32'b00010111101000010000101000101011;
		correct = 32'b10011000000000101111100001010000;
		#400 //-1.6265548 * 1.0406948e-24 = -1.6927472e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010100000010110100011101001101;
		b = 32'b11010111111000110100000001001010;
		correct = 32'b11101100011101110100011001100111;
		#400 //2392786700000.0 * -499730520000000.0 = -1.1957486e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100000110001000010011001010001;
		b = 32'b00011101111111001101001000000001;
		correct = 32'b00111111010000011011011010100000;
		#400 //1.1307259e+20 * 6.6920984e-21 = 0.7566929
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001000100010000000111011100011;
		b = 32'b11101111111010100011000110111011;
		correct = 32'b01111000111110001111000000010011;
		#400 //-278647.1 * -1.4495923e+29 = 4.0392466e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100101010000100010100101100001;
		b = 32'b00001111101000011111100000111110;
		correct = 32'b10110101011101011011000010011010;
		#400 //-5.73064e+22 * 1.5971445e-29 = -9.15266e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110000000010101110001101010;
		b = 32'b10000011011101010100110001110111;
		correct = 32'b10000001111101111110100000101010;
		#400 //0.1263291 * -7.2086806e-37 = -9.106661e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101000110100100011111011101000;
		b = 32'b11001111000011001101000011100001;
		correct = 32'b11111000011001110100101111100110;
		#400 //7.942859e+24 * -2362499300.0 = -1.8765e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000101000001111011010010111100;
		b = 32'b01110101011111010011100100101001;
		correct = 32'b11111011000001100011101111101011;
		#400 //-2171.296 * 3.2099865e+32 = -6.9698306e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010001100110011010000100110010;
		b = 32'b11001000001011100101110101010000;
		correct = 32'b01011010010100010100011100011111;
		#400 //-82479300000.0 * -178549.25 = 1.4726617e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110011100111110000111101001101;
		b = 32'b10011100101001000010100001000001;
		correct = 32'b01010000110010111111110110100000;
		#400 //-2.5204026e+31 * -1.0863015e-21 = 27379171000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111001101011011000000011001011;
		b = 32'b00110010100000011101111001111110;
		correct = 32'b11101100101100000000100101100011;
		#400 //-1.1260995e+35 * 1.5118754e-08 = -1.7025222e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100000101101100000010111001111;
		b = 32'b10100110010111101101111000010010;
		correct = 32'b10000111100111100111011011101111;
		#400 //3.0835843e-19 * -7.7322684e-16 = -2.38431e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001111101010101010100010000110;
		b = 32'b01100010000101101011000110001011;
		correct = 32'b01110010010010001110101000110011;
		#400 //5726342000.0 * 6.949512e+20 = 3.9795284e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100000010101100110100110001000;
		b = 32'b11110111010110100011010111010101;
		correct = 32'b11011000001101101100001011110100;
		#400 //1.8161422e-19 * -4.4258303e+33 = -803793730000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101010100010011110010100010111;
		b = 32'b10011011000011111110101001000001;
		correct = 32'b11000110000110110000101001001101;
		#400 //8.335234e+25 * -1.1904374e-22 = -9922.575
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110001011111000001110100001001;
		b = 32'b01110100111101111010111101000101;
		correct = 32'b11100110111100111110110010011111;
		#400 //-3.668733e-09 * 1.569888e+32 = -5.7594997e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011001110110110010100111110000;
		b = 32'b00111110101010101110110011001100;
		correct = 32'b01011001000100100101010010010011;
		#400 //7711141300000000.0 * 0.33383787 = 2574271000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011001001100110111001101001101;
		b = 32'b00110001111001000101111001110111;
		correct = 32'b11001011101000000001010011101000;
		#400 //-3156924700000000.0 * 6.6464128e-09 = -20982224.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010100001011101111010110000101;
		b = 32'b10110101011011001000111000101110;
		correct = 32'b00001010001000011010101110000010;
		#400 //-8.833175e-27 * -8.812375e-07 = 7.784125e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001011101111000000000001101111;
		b = 32'b00110101001110101101010011001000;
		correct = 32'b10000001100010010011010010010100;
		#400 //-7.241562e-32 * 6.9600037e-07 = -5.04013e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000101101011000100000000111001;
		b = 32'b11000100100010101100100100000010;
		correct = 32'b00001010101110101100001110111101;
		#400 //-1.6198394e-35 * -1110.2815 = 1.7984777e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000010010001110011011010100100;
		b = 32'b10101110111101000001011010001101;
		correct = 32'b10110001101111011111000110100001;
		#400 //49.80336 * -1.1099841e-10 = -5.528094e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001111000100100110101111100101;
		b = 32'b11100110011110100111110011101100;
		correct = 32'b00110110000011110100010011010001;
		#400 //-7.2191355e-30 * -2.95724e+23 = 2.1348717e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101100110001011011110010000010;
		b = 32'b10111101000101111111111011100001;
		correct = 32'b00101010011010101100111000011111;
		#400 //-5.6200053e-12 * -0.037108306 = 2.0854888e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101000011100001100010010110100;
		b = 32'b10110110010011000111001001100000;
		correct = 32'b00011111010000000100100001010001;
		#400 //-1.33653295e-14 * -3.0464944e-06 = 4.07174e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000000100110101100001100110010;
		b = 32'b11000000000011101001101010100100;
		correct = 32'b11000001001011000110101110000101;
		#400 //4.8363276 * -2.2281885 = -10.77625
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100101000100110000010100110101;
		b = 32'b00110000100001110001100010100110;
		correct = 32'b00010110000110110010101111001110;
		#400 //1.2751982e-16 * 9.829548e-10 = 1.2534623e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000101110101000101011000111000;
		b = 32'b11000110000101110010010010010100;
		correct = 32'b01001100011110101011101001100100;
		#400 //-6794.7773 * -9673.145 = 65726864.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101010011111000101011110101110;
		b = 32'b00010000111110011100000111110100;
		correct = 32'b10111011111101100011000001110111;
		#400 //-7.626584e+25 * 9.8512015e-29 = -0.0075131017
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101101100100110010010001111110;
		b = 32'b10001010101001111010101011000000;
		correct = 32'b00111000110000001011110111100110;
		#400 //-5.6923016e+27 * -1.6145744e-32 = 9.190645e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001010001011101100001110100110;
		b = 32'b01101111011100000110101110111001;
		correct = 32'b00111010001001000010000011110110;
		#400 //8.414593e-33 * 7.440663e+28 = 0.0006261015
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001100100010000000100110100111;
		b = 32'b01010100000101010000100110100100;
		correct = 32'b10100001000111100110010101111011;
		#400 //-2.0959927e-31 * 2560447500000.0 = -5.366679e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001101111010111110001010000110;
		b = 32'b11010100011011101110110001110001;
		correct = 32'b11100010110111000010011001110110;
		#400 //494686400.0 * -4104676200000.0 = -2.0305275e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011010001000000010010000100101;
		b = 32'b11011101111011100000101010010110;
		correct = 32'b10111000100101001110100000111010;
		#400 //3.3116422e-23 * -2.1440859e+18 = -7.1004455e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111011000001011110100110101111;
		b = 32'b00100110100101111001001110000100;
		correct = 32'b00100010000111101001010000000001;
		#400 //0.0020433476 * 1.0517714e-15 = 2.1491346e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101001011111111010110101101110;
		b = 32'b01010000001100110000001010010011;
		correct = 32'b11111010001100101100100011010110;
		#400 //-1.9318443e+25 * 12013161000.0 = -2.3207557e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111010111000000101000101011001;
		b = 32'b10100110011001010001101101100111;
		correct = 32'b01100001110010001100000011000111;
		#400 //-5.823622e+35 * -7.948747e-16 = 4.62905e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001011010001000000100101011101;
		b = 32'b10010001101100011100111011101011;
		correct = 32'b10011101100010000010100011101101;
		#400 //12847453.0 * -2.80532e-28 = -3.6041217e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011101001101111011111001000011;
		b = 32'b00010111111001101100110001101011;
		correct = 32'b10110101101001011010011110101001;
		#400 //-8.2750585e+17 * 1.4915004e-24 = -1.2342254e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011111110111101000111000101101;
		b = 32'b00000011111011110100110000001000;
		correct = 32'b00100100010100000000100011010101;
		#400 //3.207361e+19 * 1.4064613e-36 = 4.511029e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011010111001100011110110011011;
		b = 32'b00010110011011110110110100100111;
		correct = 32'b00110001110101110101010110101111;
		#400 //3.240349e+16 * 1.9340709e-25 = 6.2670646e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101001110111100111010010101111;
		b = 32'b11011000110110000010110100110110;
		correct = 32'b01000011001110111101100110111101;
		#400 //-9.879022e-14 * -1901509500000000.0 = 187.85054
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111011001001111100110011111000;
		b = 32'b11101111111001100110111101010110;
		correct = 32'b11101011100101110000101100100001;
		#400 //0.0025604349 * -1.426323e+29 = -3.652007e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100011100011001101110100011000;
		b = 32'b10011101010101001010101001101110;
		correct = 32'b01000001011010100000100110111110;
		#400 //-5.1969513e+21 * -2.8146076e-21 = 14.627378
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100101011001100001110011111111;
		b = 32'b10110000101001001100000101010000;
		correct = 32'b01010110100101000001100001010111;
		#400 //-6.791745e+22 * -1.1987513e-09 = 81416130000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011111110011011010101101111000;
		b = 32'b01001010111110010010111000100001;
		correct = 32'b00101011010010000011000011010111;
		#400 //8.710455e-20 * 8165136.5 = 7.112205e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111001000000000000001101000101;
		b = 32'b10001111001110101001101000100011;
		correct = 32'b11001000101110101001111011100111;
		#400 //4.154252e+34 * -9.200194e-30 = -382199.22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110011000110100101111101011000;
		b = 32'b00001101111011111011010100110101;
		correct = 32'b00000001100100001000110001001001;
		#400 //3.5942634e-08 * 1.4773136e-30 = 5.3098545e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101111001100010110001100001000;
		b = 32'b01110111111011011000001110010100;
		correct = 32'b01100111101001001001001111011011;
		#400 //1.6133239e-10 * 9.6347115e+33 = 1.5543911e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001000000011111110011100000000;
		b = 32'b00111010100011000010011000000001;
		correct = 32'b10000011000111011000111101100010;
		#400 //-4.3304036e-34 * 0.0010692478 = -4.630275e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011110111101001000100101010011;
		b = 32'b01111011101111000011010110010000;
		correct = 32'b11011011001100111100100000000011;
		#400 //-2.5891301e-20 * 1.9544764e+36 = -5.0603936e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110001100100110100101100100111;
		b = 32'b10111110111111101010100110100100;
		correct = 32'b00110001000100101000011000101100;
		#400 //-4.286807e-09 * -0.497388 = 2.1322064e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111111000110110011111111101;
		b = 32'b00001000000110010101001110111101;
		correct = 32'b10000000100010000011001110001001;
		#400 //-2.7108932e-05 * 4.6140197e-34 = -1.2508115e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111001000000010011000011110000;
		b = 32'b10010010011101111010001101110100;
		correct = 32'b01001011111110011111000101101001;
		#400 //-4.192493e+34 * -7.814093e-28 = 32760530.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111101110010101001010100100001;
		b = 32'b10110110000111001011011101001100;
		correct = 32'b11110100011110000000011111011010;
		#400 //3.3659797e+37 * -2.3352504e-06 = -7.8604057e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001011101001001010100110001011;
		b = 32'b00111011110110101101010000110110;
		correct = 32'b00001000000011001100000011100000;
		#400 //6.34256e-32 * 0.0066781295 = 4.235644e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101011110000011101001100101101;
		b = 32'b10101010000001101100011010100001;
		correct = 32'b00010110010011000001010111011010;
		#400 //-1.3772088e-12 * -1.1970504e-13 = 1.6485884e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000101101001110011100101001000;
		b = 32'b01100011000010011010011010011101;
		correct = 32'b10101001001100111101010011111010;
		#400 //-1.5725646e-35 * 2.5392097e+21 = -3.9930712e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000001000001101111010001111101;
		b = 32'b01011100111011100011001010100000;
		correct = 32'b11011110011110110010001111111001;
		#400 //-8.4346895 * 5.3637366e+17 = -4.5241454e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011000000011010101000101011001;
		b = 32'b11100010110101101110110100001110;
		correct = 32'b10111011011011010100100110111001;
		#400 //1.8264893e-24 * -1.9823424e+21 = -0.0036207272
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000100001001001111001101111010;
		b = 32'b01011011001110000010110111001111;
		correct = 32'b11011111111011010101100100001000;
		#400 //-659.8043 * 5.1841763e+16 = -3.420542e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101011011001111110101111010111;
		b = 32'b00010110010011100110000110100110;
		correct = 32'b01000010001110101111100000111110;
		#400 //2.8037559e+26 * 1.667136e-25 = 46.742424
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010100001110010000101100101010;
		b = 32'b00111010010010010111110100010000;
		correct = 32'b00001111000100011010010000101010;
		#400 //9.342315e-27 * 0.0007686177 = 7.180669e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100100101001011001010011011100;
		b = 32'b10111000100101010001011001000110;
		correct = 32'b01011101110000001101110000011000;
		#400 //-2.4435514e+22 * -7.1090224e-05 = 1.7371261e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000100110000110101011000110100;
		b = 32'b11010110101100101001101110011000;
		correct = 32'b01011100000010000100100010101001;
		#400 //-1562.6938 * -98190670000000.0 = 1.5344195e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001111000001111101111000001101;
		b = 32'b00111110101001111110001000000100;
		correct = 32'b10001110001100100011001110011101;
		#400 //-6.698779e-30 * 0.32789624 = -2.1965045e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010110011110110101010010111011;
		b = 32'b10010100111010110010000100010110;
		correct = 32'b10101011111001101101011101000011;
		#400 //69085333000000.0 * -2.3741986e-26 = -1.640223e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110101011101000000010100110111;
		b = 32'b11110010011100111000111110010101;
		correct = 32'b11101000011010000010100111010000;
		#400 //9.090467e-07 * -4.82422e+30 = -4.3854413e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010110000001001010110000111110;
		b = 32'b10000111101000010101101010001011;
		correct = 32'b10011110001001110011111001111111;
		#400 //36468827000000.0 * -2.4277804e-34 = -8.85383e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100001010101010011100011011110;
		b = 32'b10101101111010101011100101001011;
		correct = 32'b00001111110000111000000001001111;
		#400 //-7.224247e-19 * -2.6685007e-11 = 1.9277907e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000011101011010100111100100111;
		b = 32'b01110110110010000101100101011010;
		correct = 32'b10111011000001111010001001010100;
		#400 //-1.0186199e-36 * 2.0317805e+33 = -0.002069612
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100010110101100010101110011001;
		b = 32'b00110110100011001010110100111110;
		correct = 32'b10011001111010110110000110001110;
		#400 //-5.8050977e-18 * 4.192493e-06 = -2.4337833e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110110111110101111101110000000;
		b = 32'b10101100100100010011111001111100;
		correct = 32'b11100100000011100110010110110110;
		#400 //2.5452641e+33 * -4.128085e-12 = -1.0507067e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001100111111100100110010001010;
		b = 32'b11100100010001011010110010001001;
		correct = 32'b10110001110001000101110001001010;
		#400 //3.9180962e-31 * -1.4585764e+22 = -5.714843e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111111001101000101101110010001;
		b = 32'b00110011110110011001111010110010;
		correct = 32'b10110011100110010101000101101100;
		#400 //-0.7045222 * 1.01337164e-07 = -7.139428e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010101100011000000101111110110;
		b = 32'b01100000101100100111110001011111;
		correct = 32'b01110110110000110100100010110110;
		#400 //19247875000000.0 * 1.0289007e+20 = 1.9804153e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111100111001111101100000001000;
		b = 32'b01011111000000010011010010000000;
		correct = 32'b01011100011010100000011011010000;
		#400 //0.028301254 * 9.310207e+18 = 2.6349054e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001111000101110000101100111010;
		b = 32'b01011001011101110100111110101100;
		correct = 32'b01101001000100011110101011010111;
		#400 //2534095400.0 * 4350745000000000.0 = 1.1025203e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011001010100101000001100110110;
		b = 32'b01110011010001001100000000001101;
		correct = 32'b01001101001000011100101001100010;
		#400 //1.0883243e-23 * 1.5588157e+31 = 169649700.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100010101111100010100110001011;
		b = 32'b11110010100000010110001100010101;
		correct = 32'b11010101110000000011100100010001;
		#400 //5.154359e-18 * -5.1255487e+30 = -26418916000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001111011100111111010101000000;
		b = 32'b10111101010100100001110100001000;
		correct = 32'b01001101010010000011101011011001;
		#400 //-4092936200.0 * -0.051297218 = 209956240.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100111000010111101100000100111;
		b = 32'b10110011001101110001011100001111;
		correct = 32'b00011010110010000000100000111001;
		#400 //-1.9407301e-15 * -4.262898e-08 = 8.2731346e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100011111000011011010101110001;
		b = 32'b11001111010010000011010111101011;
		correct = 32'b10110011101100001000010101001010;
		#400 //2.4471392e-17 * -3358976800.0 = -8.219884e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001010011111101010000111011000;
		b = 32'b11000000011010100110000111100001;
		correct = 32'b10001011011010010010000101001011;
		#400 //1.22600946e-32 * -3.662224 = -4.4899215e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101100011101101011110100100011;
		b = 32'b00100100111011011100110101110011;
		correct = 32'b10010001111001010011001100011110;
		#400 //-3.5063695e-12 * 1.0313041e-16 = -3.6161333e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101111111101010100001010010101;
		b = 32'b10010000100010110011011101010111;
		correct = 32'b01000001000001010110000000101100;
		#400 //-1.5180864e+29 * -5.49111e-29 = 8.335979
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001000000001011010101101000011;
		b = 32'b01100111110000101001001010110011;
		correct = 32'b10110000010010110011000011000100;
		#400 //-4.022455e-34 * 1.8376904e+24 = -7.392027e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000011011011110000110001000100;
		b = 32'b00010010001111000111110110010000;
		correct = 32'b10010110001100000000001001000001;
		#400 //-239.04791 * 5.947711e-28 = -1.4217878e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100011011010110010001100110101;
		b = 32'b00100101000110111011101111100110;
		correct = 32'b10001001000011110000101011100111;
		#400 //-1.2746831e-17 * 1.350777e-16 = -1.7218125e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100111100111110111101000111101;
		b = 32'b10011110011000001111001101010101;
		correct = 32'b01000110100011000010001010001011;
		#400 //-1.5062223e+24 * -1.1908781e-20 = 17937.271
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110111000110101100111111111111;
		b = 32'b00000110100010000001110001100011;
		correct = 32'b10111110001001001001111101010100;
		#400 //-3.1399702e+33 * 5.1199225e-35 = -0.16076404
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101011101111010101110110000101;
		b = 32'b01000010010101111010010011110110;
		correct = 32'b11101110100111111000001110010001;
		#400 //-4.5785723e+26 * 53.911095 = -2.4683585e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111000010111111001111001010101;
		b = 32'b00011001000011010101001101111001;
		correct = 32'b10010001111101101110011000111110;
		#400 //-5.33148e-05 * 7.306386e-24 = -3.8953854e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101101101000111001110011101110;
		b = 32'b00001001011100001101111001001100;
		correct = 32'b10110111100110011111000100110010;
		#400 //-6.3294716e+27 * 2.8993473e-33 = -1.8351337e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111100010111001100110011000000;
		b = 32'b00100110101101011010111101011001;
		correct = 32'b11100011100111001011010000000000;
		#400 //-4.5858325e+36 * 1.2606926e-15 = -5.781325e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111101001100100010011110001111;
		b = 32'b11100110110000011011000101101010;
		correct = 32'b11100100100001101100101101001010;
		#400 //0.043494757 * -4.5734472e+23 = -1.9892098e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110011000000101001111100011;
		b = 32'b00111111110011101110001101111111;
		correct = 32'b00111110101101010100101011011010;
		#400 //0.21907 * 1.6163176 = 0.3540867
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001111010000111000101110100011;
		b = 32'b01101011001110001101100100101001;
		correct = 32'b11111011000011010011001000111110;
		#400 //-3280708400.0 * 2.2346786e+26 = -7.331329e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001010001100101000110101011011;
		b = 32'b01010010001000010110111000011011;
		correct = 32'b10011100111000010010111101100100;
		#400 //-8.596974e-33 * 173334250000.0 = -1.4901501e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100010010010001010100101011100;
		b = 32'b00010011000001110001011110110011;
		correct = 32'b00110101110100111100011111000110;
		#400 //9.253881e+20 * 1.705108e-27 = 1.5778867e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111101101010110010100011000101;
		b = 32'b00100111001101001010111100110001;
		correct = 32'b01100101011100011001101110011000;
		#400 //2.843871e+37 * 2.507499e-15 = 7.1310033e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000000101111011000011011011000;
		b = 32'b01010111001110001111001100010011;
		correct = 32'b01011000100010001110110011100000;
		#400 //5.9227104 * 203354140000000.0 = 1204407600000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010101111001000000111110100100;
		b = 32'b10111111000111010001000111000101;
		correct = 32'b10010101100010111110110101101100;
		#400 //9.2113143e-26 * -0.6135524 = -5.651624e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111000110111000110110100101110;
		b = 32'b00011000010111111101101001110011;
		correct = 32'b11010001110000001011111100110011;
		#400 //-3.5766242e+34 * 2.8932363e-24 = -103480190000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111110101001101000101110001010;
		b = 32'b00101000001010111110001110001011;
		correct = 32'b11100111010111111010011001111011;
		#400 //-1.1068819e+38 * 9.541747e-15 = -1.05615875e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100101100101001111000000111101;
		b = 32'b00100101100001001100110010011101;
		correct = 32'b00001011100110101000010111010100;
		#400 //2.58367e-16 * 2.3037e-16 = 5.9520004e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101001110100110000010100010011;
		b = 32'b11110101001101001011001101000001;
		correct = 32'b11011111100101001111001101010011;
		#400 //9.3711626e-14 * -2.2906473e+32 = -2.1466027e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100111000001100010010101111111;
		b = 32'b10011000001001100100100000110110;
		correct = 32'b10111111101011100100010001001110;
		#400 //6.334888e+23 * -2.1491454e-24 = -1.3614595
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011011011001010101010000100011;
		b = 32'b00100111111100110000010111000010;
		correct = 32'b01000011110110011011010000000110;
		#400 //6.455028e+16 * 6.745229e-15 = 435.40643
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011100110101111001110001001101;
		b = 32'b11101101101001011010010000010010;
		correct = 32'b01001011000010111000000111101101;
		#400 //-1.4267909e-21 * -6.407922e+27 = 9142765.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100010101001011100011101000011;
		b = 32'b11000101000101001100000100011010;
		correct = 32'b10101000010000001010100001111110;
		#400 //4.4934316e-18 * -2380.0688 = -1.0694677e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000011110010110000011100110110;
		b = 32'b11111110101001101011101001110000;
		correct = 32'b11000011000001000011101010001001;
		#400 //1.1932923e-36 * -1.1080994e+38 = -132.22865
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100011011011011110110011100111;
		b = 32'b00110100010100101110001000101110;
		correct = 32'b11011000010000111111111010001011;
		#400 //-4.388949e+21 * 1.9640058e-07 = -861992100000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111111110100101001100011101100;
		b = 32'b00011010101110101011111100011111;
		correct = 32'b10011011000110011010000001010101;
		#400 //-1.6452918 * 7.723657e-23 = -1.270767e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001000100011110011101010110001;
		b = 32'b10001011111111101010010111110011;
		correct = 32'b00010101000011100111100100010100;
		#400 //-293333.53 * -9.8086934e-32 = 2.8772185e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100000001011101010100001000101;
		b = 32'b01001110001001010100000110101011;
		correct = 32'b01101110111000010111111010000100;
		#400 //5.034154e+19 * 693136060.0 = 3.4893538e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111010001000101010101001100;
		b = 32'b11101101111100000110111000111110;
		correct = 32'b11110101101110000110010010000011;
		#400 //50261.297 * -9.3012096e+27 = -4.6749084e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110100110011010000110101001010;
		b = 32'b01011011100101111000101101010010;
		correct = 32'b01010000111100101100010011011101;
		#400 //3.8193895e-07 * 8.531181e+16 = 32583903000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110010000011010111110110010001;
		b = 32'b11100111001001110010000000100001;
		correct = 32'b11011001101110001011110101010111;
		#400 //8.235831e-09 * -7.892279e+23 = -6499947000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000111100111101111110001000011;
		b = 32'b01011000110001000011101110101011;
		correct = 32'b10100000111100111011110001100011;
		#400 //-2.3921464e-34 * 1726084400000000.0 = -4.1290465e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100101111101100001100101001111;
		b = 32'b11100011101110101110110110100110;
		correct = 32'b11001010001100111011001011011000;
		#400 //4.2691347e-16 * -6.8964375e+21 = -2944182.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110110001111001101111100000010;
		b = 32'b00100111010100010101010001111111;
		correct = 32'b11011110000110100111000001101000;
		#400 //-9.576904e+32 * 2.9050382e-15 = -2.7821273e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001111110110010001001000001001;
		b = 32'b10011001000011110101101001010001;
		correct = 32'b00101001011100110001101101010000;
		#400 //-7283675600.0 * -7.411166e-24 = 5.398053e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111101110111110011000010000001;
		b = 32'b00100101000000110101010000001110;
		correct = 32'b01100011011001001111111000110100;
		#400 //3.708371e+37 * 1.1390918e-16 = 4.224175e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001111101011000001101100001010;
		b = 32'b00001101011011000011001101011110;
		correct = 32'b10011101100111101100101101110110;
		#400 //-5774906400.0 * 7.2784946e-31 = -4.2032625e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111011111101000111100000011101;
		b = 32'b01000001011100101011101011000011;
		correct = 32'b10111101111001111100101111100101;
		#400 //-0.0074606077 * 15.170596 = -0.11318187
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000101101010101111000000011101;
		b = 32'b11001100100011111101110001111111;
		correct = 32'b11010010110000000001111010110111;
		#400 //5470.014 * -75424760.0 = -412574500000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110011010010110100101010011101;
		b = 32'b10110110000101101110101111100111;
		correct = 32'b00101001111011111011001000011010;
		#400 //-4.733248e-08 * -2.2489055e-06 = 1.0644628e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111111101000011100110111101011;
		b = 32'b00110111111101101100111100101001;
		correct = 32'b10111000000110111111111011001111;
		#400 //-1.2640966 * 2.9421952e-05 = -3.719219e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011000111100000110011011010100;
		b = 32'b01001010100111010000110110000111;
		correct = 32'b00100100000100110111101111000100;
		#400 //6.2142376e-24 * 5146307.5 = 3.1980377e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110100100111011100100100001000;
		b = 32'b01000111011011000100110011010101;
		correct = 32'b10111100100100011010010010101110;
		#400 //-2.9389798e-07 * 60492.832 = -0.01777872
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101100011011110010010100001110;
		b = 32'b00101110000110101011111100000110;
		correct = 32'b01011011000100001000111010111101;
		#400 //1.156433e+27 * 3.518521e-11 = 4.068934e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011101001001000011010110011101;
		b = 32'b00010010101001001010001100011000;
		correct = 32'b00110000010100110011010111101100;
		#400 //7.395335e+17 * 1.0390061e-27 = 7.683798e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010100100001000011111011110100;
		b = 32'b11100010110010011100101111001111;
		correct = 32'b10110111110100000111110101101101;
		#400 //1.3353424e-26 * -1.8612408e+21 = -2.4853938e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101001110101001111000100011101;
		b = 32'b11111000111010010110111001100110;
		correct = 32'b11100011010000100010101101001000;
		#400 //9.456518e-14 * -3.7876385e+34 = -3.581787e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011101100100001001000011010010;
		b = 32'b11011101110100011000001111011010;
		correct = 32'b11111011111011001010000101100001;
		#400 //1.3021321e+18 * -1.8871438e+18 = -2.4573104e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000001011101011111111100001001;
		b = 32'b10011110010010010100010011000101;
		correct = 32'b10100000010000010110011101010011;
		#400 //15.374764 * -1.0655073e-20 = -1.6381923e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101001010100000100011100000000;
		b = 32'b11100010001010001111111111100101;
		correct = 32'b01001100000010010111111011001001;
		#400 //-4.624686e-14 * -7.7937304e+20 = 36043556.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101110110101000110101110111010;
		b = 32'b11101100001100100111110000010010;
		correct = 32'b01011011100101000001100111011010;
		#400 //-9.65978e-11 * -8.630988e+26 = 8.337344e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101111000110100110111001001111;
		b = 32'b00111100011111000001000110010100;
		correct = 32'b11101100000110000000111100110000;
		#400 //-4.7794046e+28 * 0.01538505 = -7.353138e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001101100011100110100011001101;
		b = 32'b00001010000011111100001111111101;
		correct = 32'b00011000000111111111001100100010;
		#400 //298654100.0 * 6.922061e-33 = 2.067302e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011001100111110110000010011100;
		b = 32'b10101101000011011010101010100111;
		correct = 32'b10000111001100000110010011101000;
		#400 //1.6479235e-23 * -8.0528145e-12 = -1.3270422e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000001111010000111011000100001;
		b = 32'b01010011011101101110010110101100;
		correct = 32'b01010101111000000011001000010010;
		#400 //29.05768 * 1060415200000.0 = 30813207000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010000111111011010000000101000;
		b = 32'b11001101001010100110000100000111;
		correct = 32'b10011110101010001100110001111011;
		#400 //1.00037664e-28 * -178655340.0 = -1.7872263e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010000110010100110110000000001;
		b = 32'b00110001110000001011000110111011;
		correct = 32'b01000011000110000101110110001001;
		#400 //27168606000.0 * 5.608141e-09 = 152.36537
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111011111101111010010011111010;
		b = 32'b11001001101110010010110100101100;
		correct = 32'b11000110001100110010000111101011;
		#400 //0.0075575085 * -1516965.5 = -11464.4795
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100100000011001101000110001011;
		b = 32'b01110011000000001001010110110011;
		correct = 32'b01010111100011010111011000111100;
		#400 //3.053515e-17 * 1.0187534e+31 = 311077900000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011000110111001000001011101100;
		b = 32'b10101101001000000001010111011100;
		correct = 32'b00000110100010011110010010101000;
		#400 //-5.7000864e-24 * -9.099801e-12 = 5.186965e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111110101000100101000111100;
		b = 32'b10011000100100010100010000000000;
		correct = 32'b10100000111100001110110011011111;
		#400 //108692.47 * -3.7550284e-24 = -4.081433e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110111010010110000001010100110;
		b = 32'b11000100000111101111110001011100;
		correct = 32'b01111011111111000010011110000100;
		#400 //-4.117539e+33 * -635.9431 = 2.6185206e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001000100000001110110110111111;
		b = 32'b01111011011101101100110101101001;
		correct = 32'b11000100011110001001011111010010;
		#400 //-7.759614e-34 * 1.28147124e+36 = -994.3722
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011101001010111001110111000111;
		b = 32'b01011111010001100100100110101100;
		correct = 32'b11111101000001001110110101101011;
		#400 //-7.728912e+17 * 1.428814e+19 = -1.1043178e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011100111110001000100111011100;
		b = 32'b11011111100101101011110110000000;
		correct = 32'b10111101000100100101100011000001;
		#400 //1.6446899e-21 * -2.1723957e+19 = -0.035729174
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001101001100110000101101110011;
		b = 32'b11011001100101001000011010111001;
		correct = 32'b00100111010011111100000110110000;
		#400 //-5.5172415e-31 * -5225803000000000.0 = 2.883202e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011010100000100001101010010010;
		b = 32'b11010000111110101010100100111111;
		correct = 32'b11101011111111101100011111101100;
		#400 //1.831048e+16 * -33643166000.0 = -6.1602253e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110101011100010110000101000111;
		b = 32'b00111111110110110000110010111110;
		correct = 32'b10110101110011101000101000111011;
		#400 //-8.9921053e-07 * 1.7113264 = -1.5388426e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001101101110000110101011110011;
		b = 32'b11001101110101111111111010111011;
		correct = 32'b11011100000110111001100101010011;
		#400 //386752100.0 * -452974430.0 = -1.7518881e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001000000111111101000110010101;
		b = 32'b10101111001110111001010010010100;
		correct = 32'b00110111111010100011010110110011;
		#400 //-163654.33 * -1.7060336e-10 = 2.791998e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101010101010100000001011101100;
		b = 32'b00110001110011000000111110001111;
		correct = 32'b10011101000001111000010010101001;
		#400 //-3.0200094e-13 * 5.93895e-09 = -1.7935685e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011001001010110101110101001111;
		b = 32'b01010111101001101100101100101110;
		correct = 32'b11110001010111110100110100000110;
		#400 //-3014676000000000.0 * 366783160000000.0 = -1.1057324e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101001001000101110011111110100;
		b = 32'b01001101110110101101000100000010;
		correct = 32'b10110111100010110011111010000110;
		#400 //-3.6172413e-14 * 458891330.0 = -1.6599206e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000100011111011010011100100011;
		b = 32'b11000000110010110011000110010100;
		correct = 32'b10000101110010010101010010101000;
		#400 //2.9816752e-36 * -6.349802 = -1.8933047e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111101011000000011110001010010;
		b = 32'b10000110101110101101000101000000;
		correct = 32'b00000100101000111010001100011101;
		#400 //-0.054745026 * -7.027289e-35 = 3.847091e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011101111110111011001100100000;
		b = 32'b10101001101000111010101011011001;
		correct = 32'b01001000001000001110101100001000;
		#400 //-2.2671094e+18 * -7.2682915e-14 = 164780.12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100001100011010001100110111101;
		b = 32'b00110100101110000110010001011010;
		correct = 32'b11010110110010110100001110011111;
		#400 //-3.253557e+20 * 3.4345686e-07 = -111745645000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010001000010011110001101010010;
		b = 32'b01100010111100011101001101010110;
		correct = 32'b00110100100000100100000011010101;
		#400 //1.0877443e-28 * 2.2304468e+21 = 2.4261558e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000111010000001011110111010101;
		b = 32'b11110111010110100010010111100011;
		correct = 32'b10111111001001000011111000101110;
		#400 //1.4500261e-34 * -4.424567e+33 = -0.6415738
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011110100100011010001110101011;
		b = 32'b01010001000110110111001000010100;
		correct = 32'b00110000001100001101110111111110;
		#400 //1.5420164e-20 * 41727115000.0 = 6.4343897e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011001110110101011111001011010;
		b = 32'b10110011010001000001010111000010;
		correct = 32'b01001101101001111000110001010100;
		#400 //-7696355000000000.0 * -4.5654595e-08 = 351373950.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010100110011001101011100010011;
		b = 32'b01000111111110010011111100011010;
		correct = 32'b11011101010001110110111110101111;
		#400 //-7038253400000.0 * 127614.2 = -8.981811e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100010000101001000110011101110;
		b = 32'b01001100110101110110111010101101;
		correct = 32'b00101111011110100000010100101010;
		#400 //2.0132348e-18 * 112948584.0 = 2.2739202e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011101011111000011000110110101;
		b = 32'b11000000101011001111001010001100;
		correct = 32'b10011110101010100110000001010111;
		#400 //3.337762e-21 * -5.404608 = -1.8039295e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000110101101011011101000010100;
		b = 32'b00111100100000000100111101000001;
		correct = 32'b10000011101101100010101010011001;
		#400 //-6.835805e-35 * 0.015662791 = -1.07067785e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100001000111001010010101001011;
		b = 32'b11000101000111110101100100110100;
		correct = 32'b11100110110000110000001001111110;
		#400 //1.8060017e+20 * -2549.5752 = -4.6045372e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001100101001110001100001000101;
		b = 32'b10000101000101110001100110001011;
		correct = 32'b10010010010001010011111111111010;
		#400 //87605800.0 * -7.1046774e-36 = -6.2241097e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011000001111000011001010100011;
		b = 32'b10110100110011101100110101111010;
		correct = 32'b11001101100110000000011111001101;
		#400 //827702700000000.0 * -3.8519994e-07 = -318831000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000111100011010011000110001110;
		b = 32'b00110001111100001011010110100000;
		correct = 32'b10111010000001001100001010100001;
		#400 //-72291.11 * 7.0055677e-09 = -0.00050644024
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100010011001100001110001110010;
		b = 32'b11110101001010010001001100110110;
		correct = 32'b11011000000101111111101000001100;
		#400 //3.1185871e-18 * -2.1432808e+32 = -668400800000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101110010111001111111001011100;
		b = 32'b00010001011010000001000111110100;
		correct = 32'b01000000010010000101011000000011;
		#400 //1.7098551e+28 * 1.8307105e-28 = 3.1302497
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010111011010100011000011011001;
		b = 32'b00110100010111101110000001110101;
		correct = 32'b01001100010010111110001110110010;
		#400 //257495520000000.0 * 2.0757018e-07 = 53448390.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001110110110101111100111010001;
		b = 32'b00010001101100000110100100011101;
		correct = 32'b00100001000101101110010110101001;
		#400 //1836902500.0 * 2.7832685e-28 = 5.112593e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000110111000101110000101011101;
		b = 32'b11001100000101010100110110010001;
		correct = 32'b01010011100001000101000111101001;
		#400 //-29040.682 * -39138884.0 = 1136619800000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111111101001011010100100010;
		b = 32'b01101100100000101100101110010000;
		correct = 32'b11100100111110100000110100100001;
		#400 //-2.9171413e-05 * 1.2649732e+27 = -3.6901056e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011110011100110111001011111111;
		b = 32'b10101010000101001010010101111010;
		correct = 32'b00001001000011010101101111011001;
		#400 //-1.28880935e-20 * -1.3202452e-13 = 1.7015444e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100110100010111110100101001100;
		b = 32'b01000011111011001110100100001111;
		correct = 32'b11101011000000010111101001110010;
		#400 //-3.3035625e+23 * 473.82077 = -1.5652966e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101001001100001010011000011000;
		b = 32'b10010110010100010000010110110000;
		correct = 32'b01000000000100000011101110000110;
		#400 //-1.3347206e+25 * -1.688468e-25 = 2.253633
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100101001110001100111100000111;
		b = 32'b10100010011000111100011010001001;
		correct = 32'b00001000001001000110111011100110;
		#400 //-1.60296e-16 * -3.086934e-18 = 4.9482315e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000111110010111111001001101111;
		b = 32'b11011101100011111101011011011011;
		correct = 32'b10100101111001010010111100101110;
		#400 //3.0686535e-34 * -1.295589e+18 = -3.9757138e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011000011000010010110011100000;
		b = 32'b10111101011001100111001101011101;
		correct = 32'b01010110010010101011001111001010;
		#400 //-990331400000000.0 * -0.056262363 = 55718384000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100011011100001111101111101;
		b = 32'b00111110111100011110100011011011;
		correct = 32'b01000011111000010000010000111101;
		#400 //952.492 * 0.47247967 = 450.0331
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100111011000001100100001110001;
		b = 32'b01000110000010111110100010001101;
		correct = 32'b10101101111101011011001000001110;
		#400 //-3.1194904e-15 * 8954.138 = -2.7932347e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101010000011101111111110110011;
		b = 32'b11100110101011111001011011101001;
		correct = 32'b11010001010001000010101000101111;
		#400 //1.2700847e-13 * -4.1459897e+23 = -52657582000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101000111100100010111100011010;
		b = 32'b11100010111011111011111011011010;
		correct = 32'b11001100011000101100111010000110;
		#400 //2.6887824e-14 * -2.211262e+21 = -59456024.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101000110001000100001111010000;
		b = 32'b00000010010101101111101100001101;
		correct = 32'b10101011101001001101000100101000;
		#400 //-7.414678e+24 * 1.5794285e-37 = -1.1710953e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110110110001110011100000001;
		b = 32'b11111101110100100000000000100001;
		correct = 32'b11111101001100011110110110011011;
		#400 //0.42363742 * -3.4892319e+37 = -1.4781692e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101101000000011000000011111111;
		b = 32'b10101101001011110101101100001101;
		correct = 32'b01011010101100010110101001111011;
		#400 //-2.5049696e+27 * -9.967816e-12 = 2.4969074e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100001110100100111100011001100;
		b = 32'b11001101001101000101011011000101;
		correct = 32'b01101111100101000100010001000110;
		#400 //-4.8531507e+20 * -189099090.0 = 9.177264e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100001010011001010101000111001;
		b = 32'b10001100000010110100110110101110;
		correct = 32'b00101101110111101011110100001111;
		#400 //-2.359626e+20 * -1.0731546e-31 = 2.5322437e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110100000011111100010011000000;
		b = 32'b10011010100010001011011110011011;
		correct = 32'b00001111000110011000111101000101;
		#400 //-1.338949e-07 * -5.654491e-23 = 7.571075e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101101110100011010100111000110;
		b = 32'b00010100110000001101011010110011;
		correct = 32'b01000011000111011110111100101011;
		#400 //8.1109513e+27 * 1.947173e-26 = 157.93425
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000111010101001111001110111110;
		b = 32'b11101110001100110111110100110100;
		correct = 32'b01110110000101010100111010010100;
		#400 //-54515.742 * -1.3887295e+28 = 7.5707616e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111111000001101001101110110001;
		b = 32'b10101000011001001111101011100110;
		correct = 32'b11100111111100001100110100101101;
		#400 //1.7892495e+38 * -1.2710947e-14 = -2.2743056e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000010100111111101010000010110;
		b = 32'b00011100001000101000010101111000;
		correct = 32'b10011111010010101110111100010100;
		#400 //-79.91423 * 5.377381e-22 = -4.2972925e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100001110110101101101001010111;
		b = 32'b10101101111011101110010101110111;
		correct = 32'b01010000010011000011101100101000;
		#400 //-5.046404e+20 * -2.715937e-11 = 13705716000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011111011111001101010001110101;
		b = 32'b11001101000111011011010110010001;
		correct = 32'b10101101000110111100000110011101;
		#400 //5.3538816e-20 * -165370130.0 = -8.853721e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011101110100100111101011111;
		b = 32'b10010010010000110101000000000110;
		correct = 32'b00011110100011100010010010110011;
		#400 //-24420030.0 * -6.1629787e-28 = 1.5050013e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100010111100011111110101100110;
		b = 32'b00110010111001111111110101101110;
		correct = 32'b11010110010110110100101100110110;
		#400 //-2.2319623e+21 * 2.7007186e-08 = -60279020000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111111111011010010001100011110;
		b = 32'b11001001101110000011110000011000;
		correct = 32'b01001010001010101010100011101000;
		#400 //-1.8526342 * -1509251.0 = 2796090.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011111011101011010101010100011;
		b = 32'b10110101010010100001110011100110;
		correct = 32'b01010101010000011111010001100000;
		#400 //-1.770214e+19 * -7.5292917e-07 = 13328458000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011001011110111110001101000110;
		b = 32'b00101101011111101000000001011001;
		correct = 32'b11000111011110100110100111001001;
		#400 //-4431256800000000.0 * 1.4466727e-11 = -64105.785
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011011100000100110111111100011;
		b = 32'b00100101100111000100001110101000;
		correct = 32'b10000001100111110011110101001110;
		#400 //-2.1579e-22 * 2.7107532e-16 = -5.8495343e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110011011011111101100100010110;
		b = 32'b11101100011110011010100101011001;
		correct = 32'b01100000011010011110100011010000;
		#400 //-5.5843962e-08 * -1.207289e+27 = 6.74198e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101001111101000010001010000100;
		b = 32'b01011011011111010101010001011110;
		correct = 32'b01000101111100011001011010010001;
		#400 //1.0841764e-13 * 7.130593e+16 = 7730.821
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000000100000111100110010000101;
		b = 32'b01101110011001001100100101111111;
		correct = 32'b01101111011010111001001111000111;
		#400 //4.118716 * 1.7701544e+28 = 7.290763e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100001011101000111010001101100;
		b = 32'b10001010110000110001110110010011;
		correct = 32'b10101100101110100101000011101100;
		#400 //2.8183716e+20 * -1.8788942e-32 = -5.295422e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101010110010001010101111111111;
		b = 32'b00101011101111110110000101110000;
		correct = 32'b00010111000101100000010010110100;
		#400 //3.5646483e-13 * 1.3598411e-12 = 4.847355e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010111000111111011101110010110;
		b = 32'b10101101100100110100101101110011;
		correct = 32'b10000101001101111100111110010110;
		#400 //5.161244e-25 * -1.6745471e-11 = -8.642746e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001010101100101010111001001000;
		b = 32'b11001100011001111010010111010100;
		correct = 32'b00010111101000011010111100000001;
		#400 //-1.7206334e-32 * -60725070.0 = 1.0448558e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111110011011111110101101001001;
		b = 32'b10111101000000010001100100011010;
		correct = 32'b00111011111100011111101000101100;
		#400 //-0.23429598 * -0.03151808 = 0.007384559
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111000000100101011001100110010;
		b = 32'b00101111011010110011011110111000;
		correct = 32'b10101000000001101100101001101101;
		#400 //-3.4976e-05 * 2.1392921e-10 = -7.482388e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101101010001100101001011011010;
		b = 32'b11000101010110101110001001110111;
		correct = 32'b11110011001010011001000111111111;
		#400 //3.836137e+27 * -3502.154 = -1.3434743e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001001000100110001110001111000;
		b = 32'b01010011010101011000100111000111;
		correct = 32'b00011100111101010110101110111001;
		#400 //1.7707867e-33 * 917139550000.0 = 1.6240586e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010010111010111001001111100100;
		b = 32'b01011010000110011001110001011101;
		correct = 32'b10101101100011010101101101000111;
		#400 //-1.4867043e-27 * 1.0809399e+16 = -1.607038e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110001001000011101010111001001;
		b = 32'b10110001010100111100100100001111;
		correct = 32'b11100011000001011110001001001111;
		#400 //8.013686e+29 * -3.081883e-09 = -2.4697242e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101010010011110110100001111011;
		b = 32'b11011110101001000100001000111100;
		correct = 32'b01001001100001010001010010011000;
		#400 //-1.8421542e-13 * -5.9180444e+18 = 1090195.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111010100111111110000001000;
		b = 32'b01011110001000010100100101010010;
		correct = 32'b11010110000001011000111000111000;
		#400 //-1.2635261e-05 * 2.9054776e+18 = -36711468000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110010100100101100111100001100;
		b = 32'b10000001000101000111101111011111;
		correct = 32'b10110100001010100100110101111001;
		#400 //5.815695e+30 * -2.727218e-38 = -1.5860668e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110110100100010010111111101111;
		b = 32'b00001100100000000110001000111111;
		correct = 32'b01000011100100011001111101011111;
		#400 //1.4723735e+33 * 1.9780652e-31 = 291.2451
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011111010010101000011110101;
		b = 32'b00011111011001000111010100010100;
		correct = 32'b10101011110100000011011011001110;
		#400 //-30581226.0 * 4.8377723e-20 = -1.47945e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000110110000110100110111010;
		b = 32'b00101101010100110010010001011011;
		correct = 32'b10011110101100100111110111100000;
		#400 //-1.5746118e-09 * 1.2002034e-11 = -1.8898544e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000001100000000100001011001010;
		b = 32'b00010101011100111101001000000111;
		correct = 32'b00010111011101000101000101000000;
		#400 //16.032612 * 4.9239142e-26 = 7.8943204e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000110000000100110110010101000;
		b = 32'b00110011011100000010100101111010;
		correct = 32'b00111001111101001011010111111110;
		#400 //8347.164 * 5.5917077e-08 = 0.000466749
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001010110000110110001111000010;
		b = 32'b01101111100010000100100100001010;
		correct = 32'b11111010110100000000100101111100;
		#400 //-6402529.0 * 8.435652e+28 = -5.4009506e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101111111001001101010101000010;
		b = 32'b10111001100001100110011001000110;
		correct = 32'b10101001111100000100011000011000;
		#400 //4.1624487e-10 * -0.0002563467 = -1.06703004e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011011100101000110111000110001;
		b = 32'b10111110011001000111000101101010;
		correct = 32'b00011010100001000111001111100110;
		#400 //-2.4555756e-22 * -0.22308889 = 5.4781164e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010011001000011110000000010111;
		b = 32'b01010110000110010110100110101010;
		correct = 32'b01101001110000100000001101111100;
		#400 //695249340000.0 * 42169776000000.0 = 2.9318508e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111100010111111111101010111111;
		b = 32'b00101111111101001100010101011101;
		correct = 32'b01101100110101100010011110101011;
		#400 //4.6518717e+36 * 4.4523576e-10 = 2.0711796e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011101101110001101100000101011;
		b = 32'b01011000010101010011001011001111;
		correct = 32'b11110110100110011111000010001011;
		#400 //-1.6649304e+18 * 937656800000000.0 = -1.5611332e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011110100110011111011011000;
		b = 32'b00110100110100111101100000110011;
		correct = 32'b11000001001011101100111100110011;
		#400 //-27688368.0 * 3.9459118e-07 = -10.925586
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101101000000110110001111001011;
		b = 32'b01010000100000101111110110000000;
		correct = 32'b01111110000001100111010110010001;
		#400 //2.5414487e+27 * 17581212000.0 = 4.468175e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010110000101010101110100001100;
		b = 32'b11100110101100010110100011000000;
		correct = 32'b11111101010011110000010011100110;
		#400 //41056716000000.0 * -4.1889558e+23 = -1.7198477e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101010010100010001001010010100;
		b = 32'b11010011110010010101100110001001;
		correct = 32'b11111110101001000111000010110110;
		#400 //6.3188307e+25 * -1729581200000.0 = -1.0928931e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001111110101000111001100001010;
		b = 32'b00110101100011001000110001111010;
		correct = 32'b11000101111010010100011011111011;
		#400 //-7128618000.0 * 1.0471697e-06 = -7464.8726
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101001101111000011011101000100;
		b = 32'b10100000101010000111010111001101;
		correct = 32'b01001010111101111011010111000001;
		#400 //-2.844238e+25 * -2.853826e-19 = 8116960.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000110100101110011110001011010;
		b = 32'b01111100110000011000100000111111;
		correct = 32'b11000011111001001010100111111010;
		#400 //-5.6888566e-35 * 8.0390135e+36 = -457.32794
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011100111101100011011100111011;
		b = 32'b11001110110001011001100110011000;
		correct = 32'b10101100001111100000110000111010;
		#400 //1.6293191e-21 * -1657588700.0 = -2.700741e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010101110011010000001100010;
		b = 32'b01111011010101001000000101110000;
		correct = 32'b11110110100110100001011010101100;
		#400 //-0.0014162178 * 1.1033922e+36 = -1.5626437e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010011011110001111000000000011;
		b = 32'b01100000100011010110011010001101;
		correct = 32'b11110100100010010111111111101010;
		#400 //-1069178600000.0 * 8.151189e+19 = -8.715077e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110110110010111111001001100000;
		b = 32'b10101010110110101110010101111000;
		correct = 32'b01100010001011100110001100110101;
		#400 //-2.068266e+33 * -3.8883805e-13 = 8.042205e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000011110001000100001100001111;
		b = 32'b01111000100111101100100110010011;
		correct = 32'b10111100111100110111011111011001;
		#400 //-1.15352405e-36 * 2.5764729e+34 = -0.029720234
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101001000010000010111101001011;
		b = 32'b11010110101111101010001001000110;
		correct = 32'b11000000010010101101001011011010;
		#400 //3.0239086e-14 * -104802080000000.0 = -3.1691194
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011011111101101110110111101100;
		b = 32'b01101010101001011111010111110101;
		correct = 32'b01000111001000000001010010010111;
		#400 //4.085104e-22 * 1.0031713e+26 = 40980.59
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000000100000100011110011001000;
		b = 32'b01111100000010101001111001110011;
		correct = 32'b00111101000011010000101011000000;
		#400 //1.1960419e-38 * 2.8790028e+36 = 0.03443408
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100010010001110110001101100110;
		b = 32'b01001110110011000001101110010101;
		correct = 32'b10110001100111101111100010110001;
		#400 //-2.702215e-18 * 1712179800.0 = -4.626678e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110010100111010110010100110100;
		b = 32'b10011100100110101001110100110011;
		correct = 32'b10001111101111100001111100001111;
		#400 //1.8323227e-08 * -1.02315e-21 = -1.874741e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010010100100001110011001011;
		b = 32'b01100100100011010100111100101110;
		correct = 32'b11011111011001111111010110110001;
		#400 //-0.0008015155 * 2.0853571e+22 = -1.671446e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001101001010010010011010110111;
		b = 32'b11100101101110010101000010100000;
		correct = 32'b01110011011101001110010010000000;
		#400 //-177367920.0 * -1.0939063e+23 = 1.9402389e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111010100111010101011101111;
		b = 32'b10110110110001011000011100100011;
		correct = 32'b00101110101000110101001001000110;
		#400 //-1.2616379e-05 * -5.8867895e-06 = 7.4269965e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000111011000100101111011011111;
		b = 32'b11110010100101100010000110010111;
		correct = 32'b00111010100001001100000101001010;
		#400 //-1.703023e-34 * -5.94731e+30 = 0.0010128405
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100101101110001000110000010110;
		b = 32'b00101110011110101100010100111111;
		correct = 32'b01010100101101001100011011111111;
		#400 //1.08937445e+23 * 5.701861e-11 = 6211461700000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000110111101001011001101011101;
		b = 32'b00000101101000100111100001011101;
		correct = 32'b10001101000110110100110010001110;
		#400 //-31321.682 * 1.5278621e-35 = -4.785521e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111001100010001000100110101;
		b = 32'b11010000000001000110110110010101;
		correct = 32'b01000111101101110011000101010101;
		#400 //-1.0554028e-05 * -8887096000.0 = 93794.664
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101100001111011000100011100110;
		b = 32'b11110000001011000110101100100101;
		correct = 32'b11011100111111110100111010011100;
		#400 //2.693451e-12 * -2.134438e+29 = -5.749004e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111000110111100001110011010110;
		b = 32'b10111110000001011010010110111110;
		correct = 32'b11110111011001111110100110010001;
		#400 //3.6039836e+34 * -0.13051507 = -4.7037417e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000110111101001111001100000010;
		b = 32'b00010001000100001000000011101101;
		correct = 32'b10011000100010100100010000001101;
		#400 //-31353.504 * 1.1399325e-28 = -3.5740878e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100111110110011011010000100110;
		b = 32'b11100011011110101100101100111010;
		correct = 32'b11001011110101010100011011000000;
		#400 //6.0424916e-15 * -4.62633e+21 = -27954560.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000011000111101011010000011100;
		b = 32'b00110011001110001001101011001010;
		correct = 32'b10110110111001001110001011010011;
		#400 //-158.70355 * 4.298162e-08 = -6.8213353e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101100010110111000110001100010;
		b = 32'b11111011110001010111010011100011;
		correct = 32'b01101000101010010101011101000110;
		#400 //-3.11997e-12 * -2.0505065e+36 = 6.397519e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100010100110111110100011010100;
		b = 32'b00101001100011100100000011010101;
		correct = 32'b10001100101011010100010101000011;
		#400 //-4.225935e-18 * 6.3173133e-14 = -2.6696556e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110110011001000011010110111;
		b = 32'b10111110110000001100110011110010;
		correct = 32'b10111110000110100000100011000110;
		#400 //0.3994653 * -0.3765636 = -0.1504241
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100101111110000110010010100000;
		b = 32'b00010101001110110010000100100011;
		correct = 32'b10111011101101011001000110101000;
		#400 //-1.4662539e+23 * 3.779049e-26 = -0.005541045
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001100111010001111100101001100;
		b = 32'b01010010001001100000011010000110;
		correct = 32'b11011111100101110001011110010111;
		#400 //-122145380.0 * 178268500000.0 = -2.1774673e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111110010011110010010111010011;
		b = 32'b11101110111100011111010111001011;
		correct = 32'b01101101110000111100100101111111;
		#400 //-0.20229273 * -3.7441516e+28 = 7.5741463e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111101011101011110111001010001;
		b = 32'b01110011101100110111010011111010;
		correct = 32'b01110001101011000110011000000011;
		#400 //0.06004173 * 2.8436087e+31 = 1.7073519e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100000011111111010110110111101;
		b = 32'b01000001110111011110011110010011;
		correct = 32'b00100010110111011010000001000101;
		#400 //2.1656825e-19 * 27.738073 = 6.007186e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100000100001111010010100011010;
		b = 32'b10110011101000001001001101010111;
		correct = 32'b10010100101010100010101010000100;
		#400 //2.2979145e-19 * -7.4773816e-08 = -1.7182383e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111000111001100000110110111101;
		b = 32'b10011111101111110010011111101110;
		correct = 32'b10011001001010111100100000100010;
		#400 //0.000109698136 * -8.0957705e-20 = -8.880909e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110111101011100010010111010010;
		b = 32'b10101010101010010010001111101000;
		correct = 32'b01100010111001100001111011001001;
		#400 //-7.0642714e+33 * -3.0045346e-13 = 2.1224847e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110100010110101110000000101011;
		b = 32'b01110011110100101001100010110110;
		correct = 32'b11101000101101000000111001110100;
		#400 //-2.0384384e-07 * 3.3370352e+31 = -6.8023406e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000011100000000001100110000001;
		b = 32'b00110100111101010001001010101000;
		correct = 32'b00111000111101010100001101111101;
		#400 //256.19925 * 4.564838e-07 = 0.00011695081
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101100000100110101000001101011;
		b = 32'b10011010011110110011110010001101;
		correct = 32'b10000111000100001001001010110001;
		#400 //2.0934597e-12 * -5.1954496e-23 = -1.0876465e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010000110000111100101010100001;
		b = 32'b01111001100101110101001010010011;
		correct = 32'b01001010111001110111011101011001;
		#400 //7.722614e-29 * 9.821395e+34 = 7584684.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011011100111110010110011110111;
		b = 32'b00001111101110100010010000011011;
		correct = 32'b00101011111001110111101000111101;
		#400 //8.960792e+16 * 1.8354923e-29 = 1.6447465e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011110001110101100111000001101;
		b = 32'b01010101111011001001100001000100;
		correct = 32'b00110100101011001010010100010000;
		#400 //9.889368e-21 * 32517340000000.0 = 3.2157595e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110010000110010110011101001011;
		b = 32'b01000011111100111001011011011011;
		correct = 32'b00110110100100011111011101110010;
		#400 //8.929258e-09 * 487.17856 = 4.350143e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010110110001010000110011100111;
		b = 32'b11000011001011001001100101011111;
		correct = 32'b10011010100001001101101010111001;
		#400 //3.183521e-25 * -172.5991 = -5.4947286e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110110010011011110001100011110;
		b = 32'b00001010011011010101010100100101;
		correct = 32'b00000001001111101101111110111101;
		#400 //3.067958e-06 * 1.1427149e-32 = 3.5058013e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101000111111001100110100001000;
		b = 32'b01000111011011010010111101000100;
		correct = 32'b01110000111010100011100001111101;
		#400 //9.550548e+24 * 60719.266 = 5.7990226e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101001001000111011010010101111;
		b = 32'b00111101010001110111110110111100;
		correct = 32'b00100110111111110010001110110111;
		#400 //3.634999e-14 * 0.048703894 = 1.770386e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111001101011101111010101101111;
		b = 32'b10100100011000101101101110010100;
		correct = 32'b10011110100110110000101010111101;
		#400 //0.00033370728 * -4.9191928e-17 = -1.6415705e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101011111101110011100000111111;
		b = 32'b01000101010100000100101011110001;
		correct = 32'b00110001110010010010011000010010;
		#400 //1.7566017e-12 * 3332.6838 = 5.854198e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111000000110101001101011110100;
		b = 32'b11111110111110101101010101001100;
		correct = 32'b11110111100101110111110000100011;
		#400 //3.6860773e-05 * -1.6670725e+38 = -6.144958e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111011100101001010011011011110;
		b = 32'b01010101100110100010011001001101;
		correct = 32'b11010001101100110000010100111110;
		#400 //-0.0045364937 * 21186161000000.0 = -96110890000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001110001101011010101110111110;
		b = 32'b11001100011100101001110011001010;
		correct = 32'b00011011001011000010101110011110;
		#400 //-2.2392663e-30 * -63599400.0 = 1.42416e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100100110000001001101100001001;
		b = 32'b10011101011111100111111011001011;
		correct = 32'b10000010101111110111100100111000;
		#400 //8.3529367e-17 * -3.368217e-21 = -2.8134504e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101101001101000000001111111110;
		b = 32'b11011001001111000111010000101100;
		correct = 32'b11000111000001001000010010011111;
		#400 //1.0232702e-11 * -3315314200000000.0 = -33924.62
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001101010000111101111100011101;
		b = 32'b11001011000011001100000101001000;
		correct = 32'b01011000110101110110001111001100;
		#400 //-205386190.0 * -9224520.0 = 1894589000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010101001101101111101011000000;
		b = 32'b11101110111011100011111101101000;
		correct = 32'b01000100101010100100101001110001;
		#400 //-3.6952414e-26 * -3.6867043e+28 = 1362.3263
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111100110111000000011010101100;
		b = 32'b10011101100001111101110000110001;
		correct = 32'b00011010111010011000100110001001;
		#400 //-0.02685865 * -3.5961875e-21 = 9.658874e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000001010100100001000000100011;
		b = 32'b01001110101100011010001001111000;
		correct = 32'b11010000100100011100001001111001;
		#400 //-13.12894 * 1490107400.0 = -19563530000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110101000001011011000101001001;
		b = 32'b00101110110010000011001000111011;
		correct = 32'b00100100010100010001100101111001;
		#400 //4.9804345e-07 * 9.10387e-11 = 4.5341227e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001101010001100100011010011101;
		b = 32'b10111101101000011011010011101111;
		correct = 32'b10001011011110100111110100010111;
		#400 //6.109846e-31 * -0.078958385 = -4.8242356e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010101101111100111000010111111;
		b = 32'b00000010011001000100001100000101;
		correct = 32'b10011000101010011100111001000101;
		#400 //-26173931000000.0 * 1.6770028e-37 = -4.3893755e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010010010101010011110001111111;
		b = 32'b01001111000101110100011111011010;
		correct = 32'b10100001111111000000010100010001;
		#400 //-6.7285516e-28 * 2538068500.0 = -1.7077525e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101110101110010111111111011011;
		b = 32'b11001010010100110011000000001000;
		correct = 32'b11111001100110010000011100101111;
		#400 //2.8704647e+28 * -3460098.0 = -9.932089e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001000101110101111110100010011;
		b = 32'b00001101000011100011111111000111;
		correct = 32'b00010110010011111100110111101100;
		#400 //382952.6 * 4.3833898e-31 = 1.6786304e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000100000010101101000000000001;
		b = 32'b11010010010011101001101011101110;
		correct = 32'b10010110111000000000111011000110;
		#400 //1.6317333e-36 * -221840640000.0 = -3.6198475e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001000011110111010000101011011;
		b = 32'b01110010111010011001110000000010;
		correct = 32'b00111011111001011001111100110100;
		#400 //7.5722237e-34 * 9.254222e+30 = 0.007007504
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111101010001110011010011111110;
		b = 32'b00001111011010000101100110001101;
		correct = 32'b01001101001101001100110110110101;
		#400 //1.654947e+37 * 1.145573e-29 = 189586260.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101110001010001001111000110111;
		b = 32'b10100001001110000010001001001101;
		correct = 32'b10001111111100101001000010011111;
		#400 //3.83393e-11 * -6.238702e-19 = -2.3918748e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000011111000010001000101111100;
		b = 32'b01110101101101100011001000011000;
		correct = 32'b11111010001000000010111001111001;
		#400 //-450.1366 * 4.6192092e+32 = -2.0792752e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000100111010011111101101100111;
		b = 32'b10111011111011001000001101100111;
		correct = 32'b10000001010110000010101111011101;
		#400 //5.5008913e-36 * -0.007217813 = -3.9704405e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000100100110000110000000110101;
		b = 32'b10100101101110011101000011101110;
		correct = 32'b00101010110111010011001111000100;
		#400 //-1219.0065 * -3.223396e-16 = 3.9293406e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101101001101010011000011001111;
		b = 32'b00001001100001101001101111011010;
		correct = 32'b00110111001111101000101110110110;
		#400 //3.504737e+27 * 3.240589e-33 = 1.13574115e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011111110100010000110011100010;
		b = 32'b01001110100000000000001010010100;
		correct = 32'b00101110110100010001000100011000;
		#400 //8.8536256e-20 * 1073826300.0 = 9.507256e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010100111110011111001101111000;
		b = 32'b11100111101101100100010011100001;
		correct = 32'b01111101001100011111011001011000;
		#400 //-8588252700000.0 * -1.7214826e+24 = 1.4784528e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101011011110011111001111011111;
		b = 32'b01101110011000100010111000010110;
		correct = 32'b11011010010111001101011001001010;
		#400 //-8.880101e-13 * 1.7499832e+28 = -1.5540027e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001101010101011011100110000011;
		b = 32'b10101100110011000111111000001111;
		correct = 32'b10111010101010101011100100010010;
		#400 //224106540.0 * -5.812024e-12 = -0.0013025126
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000010101111101011100001000001;
		b = 32'b01100011101111101000101100111010;
		correct = 32'b00100111000011011111010001111001;
		#400 //2.8023747e-37 * 7.0298274e+21 = 1.970021e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010111100111110010001111000011;
		b = 32'b01001000000100000000100010110100;
		correct = 32'b11100000001100110001001100001101;
		#400 //-349951900000000.0 * 147490.81 = -5.1614687e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111110111011000000000000110100;
		b = 32'b11101110010111000010110110110000;
		correct = 32'b01101101110010101111101001001011;
		#400 //-0.46093905 * -1.7035484e+28 = 7.8523197e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100000100001010001011111001000;
		b = 32'b11111110001111111110001001001011;
		correct = 32'b11011111010001111000010011001000;
		#400 //2.2546814e-19 * -6.376438e+37 = -1.4376836e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101110011100010100000000110011;
		b = 32'b10011100110101010101101000001100;
		correct = 32'b00001011110010010000111101000110;
		#400 //-5.4854076e-11 * -1.4118434e-21 = 7.7445365e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001101001100000011001011110111;
		b = 32'b01101000000111011011011111101011;
		correct = 32'b11110101110110010001101110101111;
		#400 //-184758130.0 * 2.979217e+24 = -5.5043453e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001110011000100000010111100010;
		b = 32'b10011111101010010100111001110010;
		correct = 32'b00101110100101010111101100100101;
		#400 //-948009100.0 * -7.170406e-20 = 6.7976104e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010111110000110101000111010000;
		b = 32'b01011011110010111011110100100000;
		correct = 32'b00110100000110110111001000101100;
		#400 //1.2622232e-24 * 1.1469473e+17 = 1.4477035e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001111011001010111110001001000;
		b = 32'b00101100100010001101010000011110;
		correct = 32'b00111100011101010101000001011000;
		#400 //3850127400.0 * 3.8889022e-12 = 0.014972769
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011001101110001100000010111110;
		b = 32'b01010101101101110101100101111111;
		correct = 32'b10110000000001000101001001011110;
		#400 //-1.9103002e-23 * 25199376000000.0 = -4.813837e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100100010001001100010100010110;
		b = 32'b01111011011011001000000000111001;
		correct = 32'b01100000001101011100100000111111;
		#400 //4.2667663e-17 * 1.2279827e+36 = 5.2395155e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010110000011111111000011101110;
		b = 32'b11001101000100101011101001010101;
		correct = 32'b00100011101001010000000001011001;
		#400 //-1.1627472e-25 * -153855310.0 = 1.7889483e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100110000110011010000000011010;
		b = 32'b00011110001110101000110110101111;
		correct = 32'b10000100110111111110011010110010;
		#400 //-5.3299516e-16 * 9.8760575e-21 = -5.263891e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111000101101011111000110101000;
		b = 32'b10111010111101110100011011110111;
		correct = 32'b01110100001011111011111010011001;
		#400 //-2.9522097e+34 * -0.0018865754 = 5.569566e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101011110000101000010011110111;
		b = 32'b00101111110011001011101111000000;
		correct = 32'b10011100000110111001000010011110;
		#400 //-1.3821434e-12 * 3.7240788e-10 = -5.147211e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101110101001101010001111011101;
		b = 32'b10010010011000010110110001011100;
		correct = 32'b01000001100100101011110010001110;
		#400 //-2.5786305e+28 * -7.1131045e-28 = 18.342068
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111001101110000111101010010101;
		b = 32'b00000001011111000001011010001001;
		correct = 32'b10111011101101011010100011101000;
		#400 //-1.1973361e+35 * 4.6301258e-38 = -0.005543817
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000011011010101000110111101100;
		b = 32'b11101110001010000100110101100110;
		correct = 32'b10110010000110100011010000001101;
		#400 //6.892934e-37 * -1.3021763e+28 = -8.975815e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100101101011100001101101100111;
		b = 32'b11011100010101111110001110010111;
		correct = 32'b01000010100100101101001111001100;
		#400 //-3.0202757e-16 * -2.4306943e+17 = 73.413666
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011101010001011011101111101000;
		b = 32'b10110001010001100010110001011001;
		correct = 32'b11001111000110010001000110010110;
		#400 //8.905148e+17 * -2.8838e-09 = -2568066600.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010010010110100111100110000110;
		b = 32'b11010001111001010010100100101100;
		correct = 32'b11100100110000111001000111011000;
		#400 //234585420000.0 * -123029780000.0 = -2.8860994e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000111010100101110111111100111;
		b = 32'b10101011100010010110011100011100;
		correct = 32'b00110011011000100110111010110000;
		#400 //-53999.902 * -9.763054e-13 = 5.2720395e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111100100010010111000001100001;
		b = 32'b00110011110100111101001100111010;
		correct = 32'b01110000111000110111001000001101;
		#400 //5.708992e+36 * 9.863875e-08 = 5.631278e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111011010111111101010000101010;
		b = 32'b00010001010011101101100010001100;
		correct = 32'b01001101001101001101101000001111;
		#400 //1.1621854e+36 * 1.6317263e-28 = 189636850.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011100001110000101100000111110;
		b = 32'b10001001111101000101001011011010;
		correct = 32'b00100110101011111110111111000100;
		#400 //-2.0755368e+17 * -5.8818777e-33 = 1.2208053e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110001100101110000001110100011;
		b = 32'b11001010011011110100110101111011;
		correct = 32'b10111100100011010010101000011010;
		#400 //4.395092e-09 * -3920734.8 = -0.01723199
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000111100011100001110011011000;
		b = 32'b10100100010110100001101010110101;
		correct = 32'b00101100011100100010011011000111;
		#400 //-72761.69 * -4.7293836e-17 = 3.4411794e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100101011010101010011001000111;
		b = 32'b00001000011101100000000010110110;
		correct = 32'b00101110011000010111110001101111;
		#400 //6.9256315e+22 * 7.402877e-34 = 5.1269596e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010110010110100000110011010111;
		b = 32'b11000001111111110111001011101100;
		correct = 32'b11011000110110011001010010101101;
		#400 //59937170000000.0 * -31.931114 = -1913860600000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110001101101111111010111100111;
		b = 32'b00010001011010100000000100011010;
		correct = 32'b10000011101010000010011110010000;
		#400 //-5.353957e-09 * 1.8459685e-28 = -9.883236e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111011101101101011001101100100;
		b = 32'b00111000010101110111111011110110;
		correct = 32'b11110100100110011100101101000101;
		#400 //-1.897273e+36 * 5.1378236e-05 = -9.747854e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110001000010101111001111100;
		b = 32'b00111010000111101001010011110011;
		correct = 32'b10110000110001111110110001101001;
		#400 //-2.4045867e-06 * 0.0006049417 = -1.4546347e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010000101111101000011111100010;
		b = 32'b00001011010111111000011100111011;
		correct = 32'b10011100101001100101110100000011;
		#400 //-25572610000.0 * 4.3049974e-32 = -1.1009002e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010011110000110011110010110011;
		b = 32'b00101100010100101011001111100011;
		correct = 32'b11000000101000001011000011111011;
		#400 //-1677074000000.0 * 2.9942652e-12 = -5.021604
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010010100110011000110111111111;
		b = 32'b01100011011110110001101100000110;
		correct = 32'b10110110100101101001111001101111;
		#400 //-9.690662e-28 * 4.63208e+21 = -4.4887925e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110111010000001010100101101;
		b = 32'b10101100011100000100111001011111;
		correct = 32'b00100011110110011101101011100111;
		#400 //-6.916604e-06 * -3.4149556e-12 = 2.3619896e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011011111110110100011110000000;
		b = 32'b11111010101110001010110010001001;
		correct = 32'b01010111001101010100010010111111;
		#400 //-4.1570673e-22 * -4.7944103e+35 = 199306870000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110011000010110100000001010100;
		b = 32'b00111101100001110111001110001110;
		correct = 32'b10110001000100110101101110001111;
		#400 //-3.2421966e-08 * 0.06613837 = -2.144336e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100111111110101110010100010110;
		b = 32'b10100010110001000110011010101110;
		correct = 32'b10001011010000000111110000000111;
		#400 //6.9637315e-15 * -5.3234623e-18 = -3.7071163e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000100100101101101101100000010;
		b = 32'b01111011100001011001001001110110;
		correct = 32'b01000000100111010110110000101101;
		#400 //3.5465957e-36 * 1.3870921e+36 = 4.919455
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000010101001011100100010101001;
		b = 32'b10001000101010011001010011001011;
		correct = 32'b10001011110110111010001110100110;
		#400 //82.891914 * -1.0206299e-33 = -8.460196e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011100110010010100110011100110;
		b = 32'b00000011101001010100001100000111;
		correct = 32'b10100001000000011111001101000101;
		#400 //-4.5328817e+17 * 9.713217e-37 = -4.4028865e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010011101111010000011101001010;
		b = 32'b11000100000100010100101010010111;
		correct = 32'b11011000010101101001000001101001;
		#400 //1623742200000.0 * -581.16547 = -943662900000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011000010010111110000001101110;
		b = 32'b11100111011110011111010100100100;
		correct = 32'b01000000010001110001000010000101;
		#400 //-2.6350443e-24 * -1.1803913e+24 = 3.1103833
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111110101011100000000110011010;
		b = 32'b10000101001110000001011100010100;
		correct = 32'b11000100011110100100000110101101;
		#400 //1.1564699e+38 * -8.655877e-36 = -1001.0262
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000110111011010111110010100101;
		b = 32'b11001110100000001011100000110011;
		correct = 32'b01010101111011101101001001100111;
		#400 //-30398.322 * -1079777700.0 = 32823430000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001111101001111001100011000100;
		b = 32'b10011011101101001000110000001111;
		correct = 32'b00101011111011000110011000110110;
		#400 //-5623613400.0 * -2.9869013e-22 = 1.6797178e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111010010000000001100000010;
		b = 32'b00011110111110000110011010010010;
		correct = 32'b10010110110000100001001100001101;
		#400 //-1.1921629e-05 * 2.6300443e-20 = -3.1354413e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101100100101110011101101101000;
		b = 32'b00100101010101101101001010111000;
		correct = 32'b01010010011111011101000001001001;
		#400 //1.4626267e+27 * 1.8632935e-16 = 272530300000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111010100000000100100001100;
		b = 32'b00001010100111001100111101111100;
		correct = 32'b10000010011111101101110000111111;
		#400 //-1.23998725e-05 * 1.51003e-32 = -1.872418e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001010001100011101100001010110;
		b = 32'b00000101000001100000110101010010;
		correct = 32'b10001111101110100100000011111100;
		#400 //-2913813.5 * 6.303096e-36 = -1.8366047e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101111010001101010100011001011;
		b = 32'b01001110101011001111100011101100;
		correct = 32'b10111110100001100011101010010011;
		#400 //-1.8067962e-10 * 1450997200.0 = -0.26216564
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101101100011100011111111101001;
		b = 32'b01001001100011100101100000100100;
		correct = 32'b11110111100111100011000011011010;
		#400 //-5.503017e+27 * 1166084.5 = -6.416982e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110100111100101000000101110011;
		b = 32'b00011100010101001010010010101011;
		correct = 32'b00010001110010010110111100110000;
		#400 //4.51702e-07 * 7.0357744e-22 = 3.1780733e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001000100010111011000111111100;
		b = 32'b01010011110010000111100010100001;
		correct = 32'b10011100110110101100100111000000;
		#400 //-8.407602e-34 * 1722034600000.0 = -1.4478181e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010101001111001010001111000010;
		b = 32'b11101000100011101111011111110011;
		correct = 32'b00111110010100101011001100010101;
		#400 //-3.809548e-26 * -5.401199e+24 = 0.20576127
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001111010111010100100001001010;
		b = 32'b01100111000010010110010110011111;
		correct = 32'b10110110111011011000011100001101;
		#400 //-1.09100636e-29 * 6.488388e+23 = -7.0788724e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100110101011100110100100101011;
		b = 32'b11100101001001100011010100001011;
		correct = 32'b11001100011000100111100010101010;
		#400 //1.2102181e-15 * -4.9055707e+22 = -59368104.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101010010101001110110011000011;
		b = 32'b01010001111010100000010001000110;
		correct = 32'b01111100110000101010001111111000;
		#400 //6.4352587e+25 * 125636755000.0 = 8.08505e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110001001101100010000111111110;
		b = 32'b11111110101011011111110111010110;
		correct = 32'b11110000011101111001001100100001;
		#400 //2.6503808e-09 * -1.1563722e+38 = -3.0648266e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000110001110000000111100010100;
		b = 32'b01010101011111001111110101111001;
		correct = 32'b00011100001101011110010100010110;
		#400 //3.461763e-35 * 17385349000000.0 = 6.0183963e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101000001010100000101000110001;
		b = 32'b01000001101010110010111000100000;
		correct = 32'b10101010011000110110011011100100;
		#400 //-9.439106e-15 * 21.397522 = -2.0197347e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011111100000101001000101100000;
		b = 32'b01111111000001100111000000010011;
		correct = 32'b01011111000010010010001010000011;
		#400 //5.5297644e-20 * 1.7869847e+38 = 9.881605e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010100010010110011000100011000;
		b = 32'b10101101100001000111110010001010;
		correct = 32'b01000010010100100101000001010011;
		#400 //-3490808000000.0 * -1.5061969e-11 = 52.57844
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110110110010101111010100010000;
		b = 32'b10000110111100111010000101010001;
		correct = 32'b00111110010000010010011010000011;
		#400 //-2.0582313e+33 * -9.1643474e-35 = 0.18862347
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101001001100111100010000100001;
		b = 32'b10100100000110010010101001111110;
		correct = 32'b01001101110101110001110000011101;
		#400 //-1.3582745e+25 * -3.321258e-17 = 451117980.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010101110010110111110010011000;
		b = 32'b00000110101000011100010000010101;
		correct = 32'b00011101000000001001010100111000;
		#400 //27966998000000.0 * 6.0849586e-35 = 1.7017803e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000011100011000100110110011010;
		b = 32'b01011111010000001011001110100100;
		correct = 32'b01100011010100110011100101001111;
		#400 //280.60626 * 1.3885622e+19 = 3.8963925e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111100100010110011111101101111;
		b = 32'b10111010000111111000001011001010;
		correct = 32'b01110111001011011000011100010100;
		#400 //-5.784127e+36 * -0.0006084858 = 3.519559e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000100111000001001110011010111;
		b = 32'b10111101001111110010000000101000;
		correct = 32'b01000010101001111011000100111011;
		#400 //-1796.9012 * -0.046661526 = 83.84615
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011000001111010111111000100010;
		b = 32'b10101111110010101101011010101011;
		correct = 32'b10001000100101100010010001101101;
		#400 //2.4491358e-24 * -3.6896117e-10 = -9.03636e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000010000100000100000000111110;
		b = 32'b10010111100111000000010110100011;
		correct = 32'b10011010001011111101010010100110;
		#400 //36.062737 * -1.0082687e-24 = -3.6360928e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011111000100110010100101001010;
		b = 32'b00110101010011000010011011111010;
		correct = 32'b01010100111010101011011010011110;
		#400 //1.0604088e+19 * 7.605264e-07 = 8064689000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101110010101001101101101001111;
		b = 32'b11110101011101000000000010100110;
		correct = 32'b11100100010010101110000110010001;
		#400 //4.8398004e-11 * -3.0930996e+32 = -1.4969984e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101101111111110111101110100100;
		b = 32'b01000100110010010101011000011000;
		correct = 32'b00110011010010001110110111111111;
		#400 //2.9045051e-11 * 1610.6904 = 4.6782585e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111001111111000101100111100000;
		b = 32'b11101011100100100100111100010010;
		correct = 32'b11100110000100000011100100110011;
		#400 //0.00048132148 * -3.5375314e+26 = -1.7026898e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010101101110001110101000000001;
		b = 32'b00100010111011011010011111011001;
		correct = 32'b00111001001010111010100111100000;
		#400 //25414397000000.0 * 6.4416694e-18 = 0.00016371114
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111010101100100001001010001111;
		b = 32'b10011101110101011011010111001011;
		correct = 32'b10011001000101001010011111100101;
		#400 //0.0013585853 * -5.65686e-21 = -7.685327e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111111010111010011111001000111;
		b = 32'b01101010101111100101111110011001;
		correct = 32'b01101010101001001000011011010111;
		#400 //0.8642315 * 1.1507368e+26 = 9.94503e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011101101000111101111111111111;
		b = 32'b00111100101011001111100010100110;
		correct = 32'b01011010110111010111001101010101;
		#400 //1.4760546e+18 * 0.021114659 = 3.116639e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101010000111110010001101010011;
		b = 32'b00110000001101011110001001011110;
		correct = 32'b10011010111000100010000101100011;
		#400 //-1.4134292e-13 * 6.6169104e-10 = -9.352535e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101101100000100010011011011000;
		b = 32'b10111110001001000011000110011110;
		correct = 32'b10101100001001101111010000111000;
		#400 //1.4796539e-11 * -0.16034552 = -2.3725587e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111100011111011111001100011001;
		b = 32'b10011100101010101010001100111001;
		correct = 32'b11011001101010010100010101011001;
		#400 //5.274327e+36 * -1.1291848e-21 = -5955690000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101110001110100111111001011100;
		b = 32'b10011111101010111111010010110110;
		correct = 32'b00001110011110101000100101011001;
		#400 //-4.2403733e-11 * -7.282616e-20 = 3.088101e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001101011010100000110100101010;
		b = 32'b01010100011000100010001000100100;
		correct = 32'b11100010010011101011111011010110;
		#400 //-245420700.0 * 3884941600000.0 = -9.534451e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011101101111110101110001111100;
		b = 32'b11001010010100111110101001011110;
		correct = 32'b01101000100111100110100001101011;
		#400 //-1.723629e+18 * -3472023.5 = 5.9844806e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001111011010011101000110010110;
		b = 32'b11100011110110110000100001100100;
		correct = 32'b01110011110010000000110111110101;
		#400 //-3922826800.0 * -8.080883e+21 = 3.1699904e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010101010000011110110010001111;
		b = 32'b10001110100100010100010010001101;
		correct = 32'b00100100010111000001010111010101;
		#400 //-13326360000000.0 * -3.581127e-30 = 4.7723388e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100101101110100010101100010101;
		b = 32'b10100010001001110101010000101100;
		correct = 32'b10001000011100110101111010100010;
		#400 //3.229505e-16 * -2.267728e-18 = -7.3236393e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111101101100001011110101011100;
		b = 32'b00111010000101001010010111000101;
		correct = 32'b00111000010011010011111111010110;
		#400 //0.086298674 * 0.00056704535 = 4.893526e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010100101111110000111010010000;
		b = 32'b01010001010001000010011100111101;
		correct = 32'b01100110100100100110010001101111;
		#400 //6564664600000.0 * 52654494000.0 = 3.456591e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010001000110100000101110000010;
		b = 32'b00000011110010010001110001100111;
		correct = 32'b00010101011100100000100001000001;
		#400 //41351127000.0 * 1.1820239e-36 = 4.8878022e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001001100100110001101111111011;
		b = 32'b11010011100101010100110111011101;
		correct = 32'b11011101101010111001100000001111;
		#400 //1205119.4 * -1282512900000.0 = -1.5455812e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001010101001011001001101010101;
		b = 32'b11101100010100010100110100110100;
		correct = 32'b10110111100001110101111100110111;
		#400 //1.5944342e-32 * -1.0121203e+27 = -1.6137592e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100000000011101011111100110101;
		b = 32'b11001000001011110111000010001010;
		correct = 32'b01101000110000111010011011101100;
		#400 //-4.1143993e+19 * -179650.16 = 7.391525e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101000100100001000110011000011;
		b = 32'b10101100101101011011010000110110;
		correct = 32'b00010101110011010011001010001111;
		#400 //-1.6048257e-14 * -5.164337e-12 = 8.287861e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111010010000111010010111010111;
		b = 32'b01011000101111101010111111011110;
		correct = 32'b01010011100100011011101101111110;
		#400 //0.0007463372 * 1677300400000000.0 = 1251831700000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000000010000111101000111111;
		b = 32'b00011100100001011011110000001111;
		correct = 32'b10001101000011101001011110001001;
		#400 //-4.9650234e-10 * 8.849814e-22 = -4.393953e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110000110000100010110000100100;
		b = 32'b10001011001010110010011111001111;
		correct = 32'b00111100100000011101000110101110;
		#400 //-4.8074764e+29 * -3.296335e-32 = 0.015847053
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000011011100110101100110000011;
		b = 32'b11011010011011000011100001010000;
		correct = 32'b00011110011000001000110000001100;
		#400 //-7.1514036e-37 * -1.6622503e+16 = 1.1887422e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001010011111010100001000100001;
		b = 32'b11010000111000111110111001111011;
		correct = 32'b11011011111000010111110110010000;
		#400 //4149384.2 * -30592457000.0 = -1.26939854e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000011111011100101110010110;
		b = 32'b01110000010001101110010110101101;
		correct = 32'b11100001010001010010111100101001;
		#400 //-9.2330177e-10 * 2.4622277e+29 = -2.2733793e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001100100010001100101000011111;
		b = 32'b10011011010111111010100111000000;
		correct = 32'b10101000011011110000010110001010;
		#400 //71717110.0 * -1.8500977e-22 = -1.3268366e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101111011000110000111001011111;
		b = 32'b11000100100101010101011011110001;
		correct = 32'b10110100100001000111010001111010;
		#400 //2.0650635e-10 * -1194.7169 = -2.4671664e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111101110011011110011011001100;
		b = 32'b10011110101110001111010100011010;
		correct = 32'b00011101000101001100001100000101;
		#400 //-0.10053787 * -1.958313e-20 = 1.968846e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000010011111010010010000001110;
		b = 32'b10000000001110000001100010111110;
		correct = 32'b00000010110111011110000101101001;
		#400 //-63.28521 * -5.151664e-39 = 3.260241e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010010111101000001000011101011;
		b = 32'b01001110101000101010110010101100;
		correct = 32'b00100010000110110001011101010100;
		#400 //1.5402735e-27 * 1364612600.0 = 2.1018767e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110101000110001100010100001111;
		b = 32'b10101100100100100110101011111011;
		correct = 32'b11100010001011101100000001110100;
		#400 //1.9365868e+32 * -4.161447e-12 = -8.059003e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010110001100001000011010110110;
		b = 32'b10011100010010001110111110000000;
		correct = 32'b10110011000010101000111001100100;
		#400 //48523156000000.0 * -6.6483995e-22 = -3.2260132e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010000010110111000000001010111;
		b = 32'b11011011010110110101001011110010;
		correct = 32'b10101100001111000000110111101001;
		#400 //4.3289004e-29 * -6.173422e+16 = -2.6724129e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001101111010111110100000100011;
		b = 32'b01011101001001000000111111101000;
		correct = 32'b00101011100101110010111101011111;
		#400 //1.4538878e-30 * 7.3887016e+17 = 1.0742343e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011101011000001010011001100000;
		b = 32'b10111010011111000001001001010011;
		correct = 32'b10011000010111010011001111011011;
		#400 //2.9732167e-21 * -0.00096157676 = -2.858976e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111011111001010000101101101001;
		b = 32'b01000110100101001101101000101101;
		correct = 32'b11000011000001010010110111001101;
		#400 //-0.0069898856 * 19053.088 = -133.17891
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110011001010101001100010000110;
		b = 32'b00110111101001111011100100110001;
		correct = 32'b00101011010111111000100111010001;
		#400 //3.971993e-08 * 1.9994188e-05 = 7.9416774e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100010100110100110010010001000;
		b = 32'b10100100000011000101110011010000;
		correct = 32'b00000111001010010100110111101000;
		#400 //-4.1848225e-18 * -3.0436276e-17 = 1.2737041e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000110001101110011111110010011;
		b = 32'b10000111011000011000011001110000;
		correct = 32'b00001110001000010110111100011100;
		#400 //-11727.894 * -1.6966626e-34 = 1.989828e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110100100111010111101101001010;
		b = 32'b10011110000100101110000100100101;
		correct = 32'b10010011001101001011010110100001;
		#400 //2.9333233e-07 * -7.7757344e-21 = -2.2808744e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001010001101110100111010101001;
		b = 32'b01110111110111010110001101011001;
		correct = 32'b01000010100111101000011000001011;
		#400 //8.825924e-33 * 8.980567e+33 = 79.2618
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011100100010001011100101010111;
		b = 32'b11000010101100010110011010101111;
		correct = 32'b01011111101111010111110111111001;
		#400 //-3.0787504e+17 * -88.700554 = 2.7308687e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011011001101011100111110110110;
		b = 32'b00101010010001000111111001011111;
		correct = 32'b11000110000010111000110011000111;
		#400 //-5.117535e+16 * 1.7452141e-13 = -8931.194
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101100011110000101001010101000;
		b = 32'b00010100111100010100100111000100;
		correct = 32'b11000001111010100000110101011110;
		#400 //-1.20081575e+27 * 2.4363877e-26 = -29.256527
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110101000011111100111100100110;
		b = 32'b10010101010111011100000001100100;
		correct = 32'b00001010111110010010001111001111;
		#400 //-5.357309e-07 * -4.4782364e-26 = 2.3991298e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111010010101111011100101100100;
		b = 32'b00000101100110111011001101011111;
		correct = 32'b11000000100000110011010001100110;
		#400 //-2.80026e+35 * 1.464202e-35 = -4.1001463
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010100000110101100000111100010;
		b = 32'b01001100010000011100101111001111;
		correct = 32'b10100000111010100100111011000001;
		#400 //-7.81325e-27 * 50802492.0 = -3.9693257e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111011100011111000110010011110;
		b = 32'b11011101010100100101110011101001;
		correct = 32'b11011001011010111110101011100110;
		#400 //0.0043807765 * -9.473904e+17 = -4150305800000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101000001011111110100000011101;
		b = 32'b01000111011000110011110100100111;
		correct = 32'b00110000000111000010010011010111;
		#400 //9.764783e-15 * 58173.152 = 5.680482e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011110010100110111110110001010;
		b = 32'b10010001000100101101111011111000;
		correct = 32'b00101111111100101010101110011001;
		#400 //-3.809872e+18 * -1.1586077e-28 = 4.414147e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110010110011111011101000111011;
		b = 32'b00000011000111101001101110111011;
		correct = 32'b00110110100000001011001101001110;
		#400 //8.2289326e+30 * 4.6610797e-37 = 3.835571e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011010010010101100101110111111;
		b = 32'b01000000111010110111011101101011;
		correct = 32'b00011011101110101000011110100010;
		#400 //4.1937206e-23 * 7.3583274 = 3.085877e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111011100100111010010110000010;
		b = 32'b10111100001000010001010000001110;
		correct = 32'b00111000001110011100110101010000;
		#400 //-0.004505814 * -0.009831442 = 4.429865e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111100011000110000101101110;
		b = 32'b01011001110001110011011000000100;
		correct = 32'b11010001110110100111101010110111;
		#400 //-1.673467e-05 * 7009114000000000.0 = -117295210000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101010111110000111101111011001;
		b = 32'b00000111011101100100001010001111;
		correct = 32'b00110010111011110000011110011101;
		#400 //1.5019923e+26 * 1.8526543e-34 = 2.7826724e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001000001011000100001101001011;
		b = 32'b11001111011010111001010011010100;
		correct = 32'b00011000000111101000010111101011;
		#400 //-5.183847e-34 * -3952399400.0 = 2.0488633e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011011100001001110110011000111;
		b = 32'b11001111000010000001101100010101;
		correct = 32'b11101011000011010101011110110011;
		#400 //7.483007e+16 * -2283476200.0 = -1.7087269e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000010110111110010010110010000;
		b = 32'b10010111001001111000000100000001;
		correct = 32'b00011010100100100000000111110100;
		#400 //-111.573364 * -5.4123436e-25 = 6.038734e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010001011000001110110110001010;
		b = 32'b10011000010111100100111111011011;
		correct = 32'b10101010010000110101010000100111;
		#400 //60378620000.0 * -2.8733144e-24 = -1.7348675e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001010011010100111010010001011;
		b = 32'b01000110011000010000101000000001;
		correct = 32'b01010001010011100001100110011000;
		#400 //3841314.8 * 14402.501 = 55324540000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000100000010000010111011011000;
		b = 32'b11000011000011101100010011100100;
		correct = 32'b00000111100101111110010101110010;
		#400 //-1.6008233e-36 * -142.7691 = 2.285481e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001001000000101011111001001001;
		b = 32'b01100100100000101000101000001000;
		correct = 32'b10101110000001010101011000111111;
		#400 //-1.5737652e-33 * 1.9264183e+22 = -3.03173e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100010001000110111010100100111;
		b = 32'b01111100100011011100111000000011;
		correct = 32'b11011111001101010001011000100001;
		#400 //-2.215264e-18 * 5.890338e+36 = -1.3048653e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000111000111000010010110000101;
		b = 32'b11100100101110000101010111010110;
		correct = 32'b01101100011000001101111010100101;
		#400 //-39973.52 * -2.7203088e+22 = 1.0874032e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001100001101111000110111011000;
		b = 32'b01010001001111110000110111101001;
		correct = 32'b10011110000010001111110011001101;
		#400 //-1.4140492e-31 * 51285758000.0 = -7.252058e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011110000011001001011111110100;
		b = 32'b00111010011100011100101100100100;
		correct = 32'b11011001000001001100101010011101;
		#400 //-2.5327085e+18 * 0.0009223691 = -2336092000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101000011000110000101110110110;
		b = 32'b11110111111111101010101111010110;
		correct = 32'b01100000111000011101111000000101;
		#400 //-1.2603571e-14 * -1.03306926e+34 = 1.3020361e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011101011011000010000111000111;
		b = 32'b11111001110011001101110000011010;
		correct = 32'b11010111101111001111010111110000;
		#400 //3.1251802e-21 * -1.3296159e+35 = -415528960000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101000111000010111010101010111;
		b = 32'b10010000111110111011000110010110;
		correct = 32'b00111010010111011010101001110011;
		#400 //-8.517576e+24 * -9.927566e-29 = 0.000845588
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010111001000110001011010110100;
		b = 32'b00110010100011010100100000111111;
		correct = 32'b01001010001101000000001100001111;
		#400 //179317900000000.0 * 1.6447414e-08 = 2949315.8
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011011111010010010110111101110;
		b = 32'b01101011011111011100100010111100;
		correct = 32'b01000111111001110010100100111011;
		#400 //3.8576298e-22 * 3.0680617e+26 = 118354.46
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011100001010110000001000000101;
		b = 32'b01011001111111001011111100000010;
		correct = 32'b10110110101010001101010110010101;
		#400 //-5.6581764e-22 * 8892713700000000.0 = -5.0316544e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100000011111011011001101111101;
		b = 32'b10110000000110101110100010001111;
		correct = 32'b00010001000110011000010001110010;
		#400 //-2.1489321e-19 * -5.635536e-10 = 1.2110385e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001110000011001111010111011001;
		b = 32'b01101111100000100000101100101001;
		correct = 32'b01111110000011110011010111111011;
		#400 //591230500.0 * 8.049309e+28 = 4.758997e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111111111100011000000110001011;
		b = 32'b00110010001010011111101111001110;
		correct = 32'b10110010101000000101110000010001;
		#400 //-1.8867658 * 9.8943485e-09 = -1.8668318e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101001001010110110010101100011;
		b = 32'b01101111001010011110001000111110;
		correct = 32'b01011000111000110111101011001111;
		#400 //3.8057566e-14 * 5.2576477e+28 = 2000932800000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100011010010010110101100011010;
		b = 32'b10001100011100000100100010100100;
		correct = 32'b10110000001111010000110110010000;
		#400 //3.715513e+21 * -1.8510787e-31 = -6.8777073e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011011010010011011110111100010;
		b = 32'b01000100101101110110001100011011;
		correct = 32'b11100000100100001000010011010110;
		#400 //-5.678525e+16 * 1467.097 = -8.330947e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101011111010110101011000100110;
		b = 32'b01001011011101001100001001001011;
		correct = 32'b01110111111000010000000010111000;
		#400 //5.690088e+26 * 16040523.0 = 9.127198e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001110110110011111101100110000;
		b = 32'b10010011110011100100111110001100;
		correct = 32'b00100011001011111010101111011100;
		#400 //-1828558800.0 * -5.208015e-27 = 9.523162e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100110011000101110111011011101;
		b = 32'b01010101011011110001111100101100;
		correct = 32'b10111100010100111111100010100010;
		#400 //-7.873322e-16 * 16432323000000.0 = -0.012937697
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001100101000011100101101000110;
		b = 32'b01000000011010010101110000001001;
		correct = 32'b00001101100100110111110000101101;
		#400 //2.4928318e-31 * 3.6462424 = 9.089469e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110101100101111111001101110111;
		b = 32'b10000110010001110001011010101010;
		correct = 32'b00111100011011000101011101101011;
		#400 //-3.8524164e+32 * -3.744439e-35 = 0.014425139
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000010010100001000010111101010;
		b = 32'b00000101110010100111111110111101;
		correct = 32'b00001000101001001111000110110111;
		#400 //52.130775 * 1.9042912e-35 = 9.927218e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000101100101000100101011010001;
		b = 32'b01110001011110101100001111110010;
		correct = 32'b01110111100100010100001010010001;
		#400 //4745.352 * 1.2417302e+30 = 5.8924467e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101111000101001010000011000010;
		b = 32'b00011101111111110101000000111101;
		correct = 32'b00001101100101000011101010110111;
		#400 //1.3517634e-10 * 6.7580902e-21 = 9.135339e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101110110110001010000100111100;
		b = 32'b10101011001111100101100010111001;
		correct = 32'b10011010101000010001001010111111;
		#400 //9.851184e-11 * -6.762469e-13 = -6.6618325e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011100011001010010011111011101;
		b = 32'b10111101011001100001100010111111;
		correct = 32'b11011010010011011111011111110111;
		#400 //2.580064e+17 * -0.056175943 = -1.4493753e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100011101001111110011110011000;
		b = 32'b11110010100011100011100011111110;
		correct = 32'b11010110101110101000111110101111;
		#400 //1.820426e-17 * -5.6340187e+30 = -102563140000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110011010111101000000001010;
		b = 32'b00101001010110001111010111100100;
		correct = 32'b00101000010001111101101000001001;
		#400 //0.2302858 * 4.817491e-14 = 1.1093998e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101101100101001100001110100100;
		b = 32'b00100011101111001000011100110000;
		correct = 32'b10010001110110110001110001110111;
		#400 //-1.6912534e-11 * 2.0440255e-17 = -3.456965e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000001000010011010100010000010;
		b = 32'b01000000000110100010110111000110;
		correct = 32'b10000001101001011100111111110111;
		#400 //-2.5283824e-38 * 2.4090438 = -6.090984e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010000010010010100010101011011;
		b = 32'b10010010000011100011011101110001;
		correct = 32'b00100010110111111010000000011110;
		#400 //-13507063000.0 * -4.4875636e-28 = 6.06138e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001110100100100000001111010110;
		b = 32'b10011100110111101100101000101100;
		correct = 32'b10101011111111100010010101000111;
		#400 //1224862500.0 * -1.4742988e-21 = -1.8058132e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000110011110101111101001001010;
		b = 32'b11101000001100000001110101100000;
		correct = 32'b00101111001011001010100011011111;
		#400 //-4.7203657e-35 * -3.3267135e+24 = 1.5703304e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101001000001100010000100011000;
		b = 32'b10100101101000100010111000100111;
		correct = 32'b00001111001010011111001000111111;
		#400 //-2.978268e-14 * -2.8133794e-16 = 8.378998e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011100111101010111000111011000;
		b = 32'b01010110101010110011001101100111;
		correct = 32'b01110100001001000010010001010100;
		#400 //5.5269233e+17 * 94118630000000.0 = 5.2018647e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011101111110011010011000100011;
		b = 32'b01011101000101011011101100011001;
		correct = 32'b01111011100100100000010000100111;
		#400 //2.248638e+18 * 6.743278e+17 = 1.5163191e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001111011010110010110010111001;
		b = 32'b10000100000001001110000001111101;
		correct = 32'b00010011111101000010001010010011;
		#400 //-3945576700.0 * -1.5619605e-36 = 6.1628352e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101011011011010101010001101110;
		b = 32'b00111010000000111111101101000101;
		correct = 32'b00100101111101001011011001001100;
		#400 //8.4316484e-13 * 0.00050346955 = 4.2450782e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010101101111111001101010101111;
		b = 32'b11000010010100101010000000100001;
		correct = 32'b11011000100111011010010010111101;
		#400 //26333885000000.0 * -52.656376 = -1386647000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000101011011100100001011011110;
		b = 32'b11100101111110010100100110010001;
		correct = 32'b01101011111010000000001110000010;
		#400 //-3812.1792 * -1.4715329e+23 = 5.609747e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000010011000000001000000001110;
		b = 32'b10100011110000000100001001101110;
		correct = 32'b00100110101010000100011000101111;
		#400 //-56.01568 * -2.0844816e-17 = 1.1676365e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110110110000000100101001110100;
		b = 32'b00010001010101101110001011101011;
		correct = 32'b11001000101000010110100010101111;
		#400 //-1.9500607e+33 * 1.6951548e-28 = -330565.47
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011010101111010011000111000010;
		b = 32'b10101111000111100001100010100101;
		correct = 32'b10001010011010011010110111011001;
		#400 //7.8248956e-23 * -1.4378772e-10 = -1.1251239e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001101111101101111101110001000;
		b = 32'b01001110110000111101001100111001;
		correct = 32'b10011101001111001110110101100001;
		#400 //-1.5221474e-30 * 1642699900.0 = -2.5004315e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010011110111111100111001000110;
		b = 32'b01001001001101101010001101101001;
		correct = 32'b01011101100111111010101110000010;
		#400 //1922476800000.0 * 748086.56 = 1.4381791e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100000111000110010011010100110;
		b = 32'b01100100110100101110000000001010;
		correct = 32'b01000110001110110001110001111111;
		#400 //3.848087e-19 * 3.111968e+22 = 11975.124
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011011001111110000000000010011;
		b = 32'b00110000011110011001011010101001;
		correct = 32'b10001100001110100011011101111011;
		#400 //-1.5799174e-22 * 9.0799773e-10 = -1.4345614e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110000111010001010110000000110;
		b = 32'b01000010011100010100001111111110;
		correct = 32'b01110011110110110100011110111110;
		#400 //5.760679e+29 * 60.3164 = 3.4746341e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111000111000100101000010011101;
		b = 32'b11001100011011101001111101000111;
		correct = 32'b01000101110100101111001111000001;
		#400 //-0.00010791535 * -62553372.0 = 6750.469
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001111110110010011001001001100;
		b = 32'b10011011011101011101000010100010;
		correct = 32'b10101011110100001000111000100101;
		#400 //7287904000.0 * -2.0333338e-22 = -1.4818742e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110011111010111100101111011011;
		b = 32'b10111011100010101001101010100001;
		correct = 32'b01101111111111110101010010100010;
		#400 //-3.7363417e+31 * -0.004229859 = 1.5804198e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011110011010010101011101100100;
		b = 32'b10100011101000101011101001110111;
		correct = 32'b01000010100101000101001101000011;
		#400 //-4.2035044e+18 * -1.7643046e-17 = 74.16262
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111100000000010110000000011100;
		b = 32'b00001110110101000101010110000100;
		correct = 32'b11001011010101101001110110011110;
		#400 //-2.6870225e+36 * 5.2344384e-30 = -14065054.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011010100110111111000101101111;
		b = 32'b01100011011101101001110100011000;
		correct = 32'b11111110100101100011100110110010;
		#400 //-2.194704e+16 * 4.5492188e+21 = -9.984189e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111000011100011100010100111111;
		b = 32'b00110011010100011001110001000011;
		correct = 32'b01101100010001011111010110011100;
		#400 //1.9614753e+34 * 4.8803724e-08 = 9.57273e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110111010011000011000100010000;
		b = 32'b10110001111111110000000101110011;
		correct = 32'b01101001110010110110011000000111;
		#400 //-4.1414987e+33 * -7.4216415e-09 = 3.073672e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011101110010010010110101010010;
		b = 32'b00101100110110011010010100010010;
		correct = 32'b10001011001010110000100100100011;
		#400 //-5.3251117e-21 * 6.1858374e-12 = -3.2940276e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100100001011011000001010000010;
		b = 32'b00101100000001110111110110111000;
		correct = 32'b10010000101101111010101000010000;
		#400 //-3.762394e-17 * 1.9254442e-12 = -7.2442796e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010100001101001110001010001111;
		b = 32'b00010101100001100001001001101100;
		correct = 32'b00101010001111010111011100110110;
		#400 //3107580500000.0 * 5.4151234e-26 = 1.6827932e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110010101001110100001010111111;
		b = 32'b10110010111101100111000011110100;
		correct = 32'b10100110001000010000001111110000;
		#400 //1.9471711e-08 * -2.8689534e-08 = -5.586343e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100001100111001110110000110100;
		b = 32'b10101000000100100011111000010100;
		correct = 32'b01001010001100110100100110000110;
		#400 //-3.6183904e+20 * -8.118089e-15 = 2937441.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110110001100001101011100101100;
		b = 32'b10001011010000000110111010010101;
		correct = 32'b01000010000001001110110111000100;
		#400 //-8.9668794e+32 * -3.7061048e-32 = 33.232193
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111001110010110111111001000001;
		b = 32'b00110101110110100010111001111110;
		correct = 32'b01110000001011010110111001111000;
		#400 //1.3207462e+35 * 1.6255797e-06 = 2.1469782e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010001100001110000101001001110;
		b = 32'b01100101100001111100011110110110;
		correct = 32'b01110111100011110011111110010000;
		#400 //72499180000.0 * 8.015044e+22 = 5.810841e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110100011001100011111100110111;
		b = 32'b00100101011000000110101111110101;
		correct = 32'b10011010010010011101100001101001;
		#400 //-2.1443417e-07 * 1.946548e-16 = -4.174064e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110101100110010100111000100110;
		b = 32'b10101111011111000010101100111100;
		correct = 32'b00100101100101110000001011010001;
		#400 //-1.1422133e-06 * -2.2934626e-10 = 2.6196233e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111101000000011011011001110000;
		b = 32'b01100001100101100101010000011011;
		correct = 32'b01011111000110000101011100000110;
		#400 //0.031668127 * 3.46634e+20 = 1.0977249e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011001001011001010001000101100;
		b = 32'b01100011001011001100111110001100;
		correct = 32'b01111100111010010001000111010110;
		#400 //3037000400000000.0 * 3.1877953e+21 = 9.6813354e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110010011011001100101011011100;
		b = 32'b01011010011000110110101101100010;
		correct = 32'b11001101010100100101101100110101;
		#400 //-1.3783133e-08 * 1.6003222e+16 = -220574540.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000001010101000100001101111010;
		b = 32'b01010010010001101001110000111110;
		correct = 32'b00010100001001001010110110111101;
		#400 //3.8986662e-38 * 213256210000.0 = 8.314148e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100010111110101100000010011100;
		b = 32'b00010100001101001001100110000011;
		correct = 32'b00110111101100001110010111001011;
		#400 //2.3127825e+21 * 9.1179525e-27 = 2.108784e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011110110110011111001011111001;
		b = 32'b10110010000010011001011101000011;
		correct = 32'b10010001011010100100011110011101;
		#400 //2.307626e-20 * -8.0088425e-09 = -1.8481413e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001001001010001110010101101011;
		b = 32'b11011100100101010010101011010000;
		correct = 32'b01100110010001001101001110001100;
		#400 //-691798.7 * -3.3589475e+17 = 2.3237155e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100000100011100100100011101011;
		b = 32'b10010001001010110010100111101000;
		correct = 32'b10110010001111100100001111111111;
		#400 //8.202162e+19 * -1.3502435e-28 = -1.1074916e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111100011001111010001011011000;
		b = 32'b01011001001001001000101001000110;
		correct = 32'b01010110000101001110000101101111;
		#400 //0.014137946 * 2894620600000000.0 = 40923988000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101101001001000111110101101011;
		b = 32'b10111000010000111010110100111110;
		correct = 32'b01100101111110110111010110110010;
		#400 //-3.1816977e+27 * -4.6652967e-05 = 1.48435635e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000101001111111011100001110011;
		b = 32'b01000011101010111010110001011111;
		correct = 32'b10001001100000001001000101001100;
		#400 //-9.014655e-36 * 343.34665 = -3.0951516e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111101001000011101001000010011;
		b = 32'b10100111011001100101110010100011;
		correct = 32'b10100101000100011001110101001100;
		#400 //0.039506983 * -3.196913e-15 = -1.263004e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101010110010001001000110010001;
		b = 32'b01010101000011011101100110001101;
		correct = 32'b11000000010111100100010100111101;
		#400 //-3.5628144e-13 * 9747845000000.0 = -3.472976
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011101111110110010000100110100;
		b = 32'b11010110111110010000111000111110;
		correct = 32'b01110101011101000101000101000100;
		#400 //-2.2619752e+18 * -136919780000000.0 = 3.0970915e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001010011100100011101001001001;
		b = 32'b10010111000011001101111001110111;
		correct = 32'b10100010000001010100101001011111;
		#400 //3968658.2 * -4.551723e-25 = -1.8064233e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000011001111100101001110010001;
		b = 32'b10101110101110010101100111001110;
		correct = 32'b00110010100010011100110100101000;
		#400 //-190.32643 * -8.4287785e-11 = 1.6042193e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000000010011010001101011110101;
		b = 32'b01001100111110110011010000011000;
		correct = 32'b10001101100101110101001000111110;
		#400 //-7.081004e-39 * 131702980.0 = -9.325893e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011110001010000010001101001101;
		b = 32'b11011101010110010100001001011011;
		correct = 32'b11111100000011101011000110000001;
		#400 //3.028903e+18 * -9.7844846e+17 = -2.9636254e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011111110101100111101010001000;
		b = 32'b10000001010110000101010000000000;
		correct = 32'b00100001101101010011110111000011;
		#400 //-3.090963e+19 * -3.97332e-38 = 1.2281385e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001101001011001000000010011111;
		b = 32'b11100001100011011010111001110100;
		correct = 32'b11101111001111101111000011001010;
		#400 //180881900.0 * -3.266952e+20 = -5.909325e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001110110010011000011100000011;
		b = 32'b10111100011100011101111000111100;
		correct = 32'b11001011101111100110011100001100;
		#400 //1690534300.0 * -0.014762457 = -24956440.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111101010000010000001101101100;
		b = 32'b11101100010101110000110101110001;
		correct = 32'b01101010001000100010010000000010;
		#400 //-0.047122404 * -1.0399301e+27 = 4.9004006e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111001010111010001111001000101;
		b = 32'b00010111010001001000100100000110;
		correct = 32'b01010001001010011100000110000111;
		#400 //7.175697e+34 * 6.3503964e-25 = 45568520000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001110001110011000011010000010;
		b = 32'b00010100010010111110101001111110;
		correct = 32'b00100011000100111100011110011001;
		#400 //778150000.0 * 1.0295126e-26 = 8.0111524e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100101000110011101100011110110;
		b = 32'b11010100010101111101101100001111;
		correct = 32'b11111010000000011011100011011100;
		#400 //4.540777e+22 * -3708372600000.0 = -1.6838892e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111000010010100101000001111100;
		b = 32'b10101000011000111011010011010100;
		correct = 32'b11100001001100111111010001000110;
		#400 //1.6413693e+34 * -1.2640242e-14 = -2.0747306e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110001011100010011101000111111;
		b = 32'b10110110010011011110111011101010;
		correct = 32'b00101000010000100000110011000101;
		#400 //-3.5103225e-09 * -3.0686447e-06 = 1.0771932e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100101101101010110010101110001;
		b = 32'b00010010011010110101110111010011;
		correct = 32'b10111000101001101100011010011010;
		#400 //-1.0707745e+23 * 7.426857e-28 = -7.952489e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100110111001100100100111110111;
		b = 32'b11010100111000100011101111100111;
		correct = 32'b10111100010010111000001100101111;
		#400 //1.5979504e-15 * -7773341000000.0 = -0.012421413
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011100111001101000011101101101;
		b = 32'b10011011110001001110110110011111;
		correct = 32'b00111001001100010101010110101010;
		#400 //-5.1910517e+17 * -3.257904e-22 = 0.00016911948
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111100100111111011100110000101;
		b = 32'b00010111101101010110101100111111;
		correct = 32'b00010100111000100110001000101010;
		#400 //0.019497642 * 1.1723924e-24 = 2.2858887e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000110001110000010100001110001;
		b = 32'b10111011000100101101100110001010;
		correct = 32'b11000001110100110100011100011100;
		#400 //11786.11 * -0.0022407495 = -26.409721
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011111000001100111100001100100;
		b = 32'b00011110000100011111010010101110;
		correct = 32'b00111101100110010101010101101110;
		#400 //9.689605e+18 * 7.726835e-21 = 0.074869975
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100110101110000010011011010110;
		b = 32'b01110111010111000100010011010101;
		correct = 32'b01011110100111100111001011100011;
		#400 //1.2778091e-15 * 4.4675835e+33 = 5.708719e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110011110100101000100101010101;
		b = 32'b00101010001010101010100001101111;
		correct = 32'b00011110100011000101100110111000;
		#400 //9.8038676e-08 * 1.515747e-13 = 1.4860183e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100110111111100010011010110101;
		b = 32'b11010110101101010111100010110111;
		correct = 32'b10111110001101000010100100110110;
		#400 //1.7635282e-15 * -99765035000000.0 = -0.17593846
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100000001000110111010100000010;
		b = 32'b00100110101001011010011111010111;
		correct = 32'b10000111010100111000101100101010;
		#400 //-1.3845352e-19 * 1.1494668e-15 = -1.5914772e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100010100010111000011110110101;
		b = 32'b10100010000100100000000110001010;
		correct = 32'b00000101000111110010100001111000;
		#400 //-3.781971e-18 * -1.9787504e-18 = 7.483577e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001110101111010101001100111111;
		b = 32'b01110010100101110001111000100111;
		correct = 32'b01000001110111111000010011001110;
		#400 //4.667226e-30 * 5.986392e+30 = 27.939846
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010110010001001000110001010011;
		b = 32'b10000001000110010111111111100001;
		correct = 32'b10010111111010111011010000011000;
		#400 //54026740000000.0 * -2.819341e-38 = -1.5231981e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000110101101000110011011101010;
		b = 32'b01011110101001100010001001001101;
		correct = 32'b00100101111010100010010111001111;
		#400 //6.7859693e-35 * 5.9856077e+18 = 4.061815e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101010011000010001001100111100;
		b = 32'b00101010101001110110011101010111;
		correct = 32'b10010101100100110010111001100111;
		#400 //-1.9990688e-13 * 2.9736866e-13 = -5.944604e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011000000000011110011111110010;
		b = 32'b10101111000100001100111000010000;
		correct = 32'b11000111100100101111011000010010;
		#400 //571332800000000.0 * -1.3169932e-10 = -75244.14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100000111111100111111010100010;
		b = 32'b10111010011101010101101110011010;
		correct = 32'b11011011111100111110101001000001;
		#400 //1.4670618e+20 * -0.0009359658 = -1.3731197e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010001101010111001110001000100;
		b = 32'b01101000110011111101111101001100;
		correct = 32'b00111011000010110101100100001011;
		#400 //2.707535e-28 * 7.8531917e+24 = 0.002126279
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010000011110011110111101111000;
		b = 32'b00101000010010000010010101000000;
		correct = 32'b10111001010000110110011101110100;
		#400 //-16772882000.0 * 1.11103076e-14 = -0.00018635188
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101100010001101100110100000011;
		b = 32'b10011000101100010110111010001101;
		correct = 32'b10000101100010011100100110011001;
		#400 //2.8251297e-12 * -4.5865055e-24 = -1.2957473e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011011111001111100110101100010;
		b = 32'b11010110011011100110100110011001;
		correct = 32'b11110010110101111110000010001111;
		#400 //1.3049308e+17 * -65534326000000.0 = -8.551776e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011001100110100111010010110001;
		b = 32'b11101110111100111110011011101000;
		correct = 32'b11001001000100110010100000010101;
		#400 //1.5970358e-23 * -3.7742003e+28 = -602753.3
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000110111001011011010110001100;
		b = 32'b10111001101101110000110110101000;
		correct = 32'b00000001001001000100000100001000;
		#400 //-8.6406985e-35 * -0.00034914655 = 3.01687e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111010001111111110110001001101;
		b = 32'b10000000010001001110100110011000;
		correct = 32'b00111010110011101010011110010010;
		#400 //-2.4913036e+35 * -6.328611e-39 = 0.0015766493
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010011010000101101010101011110;
		b = 32'b01111110110100010001001000101101;
		correct = 32'b01010010100111110001111000000111;
		#400 //2.459144e-27 * 1.3895151e+38 = 341701800000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010011010100101101101101101010;
		b = 32'b00000111110000011110110010010100;
		correct = 32'b10011011100111111011101001000111;
		#400 //-905624300000.0 * 2.917846e-34 = -2.6424722e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011100110101111101101101110110;
		b = 32'b11010111111001111000100001011001;
		correct = 32'b10110101010000110011100111111111;
		#400 //1.4284236e-21 * -509145600000000.0 = -7.2727556e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001100001011001001111010100110;
		b = 32'b01000010001101101000110011101111;
		correct = 32'b10001110111101100010111110100100;
		#400 //-1.329814e-31 * 45.63763 = -6.068956e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001001011000110101010010110110;
		b = 32'b11101100110011100110110111000111;
		correct = 32'b10110110101101110100111110100110;
		#400 //2.7363962e-33 * -1.996457e+27 = -5.4630973e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000101100101000001011110101000;
		b = 32'b11011111001111010101011110111100;
		correct = 32'b00100101010110110001000001110000;
		#400 //-1.3926543e-35 * -1.364358e+19 = 1.9000791e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101000000110001011001110101010;
		b = 32'b10110001011001010110001011000101;
		correct = 32'b00011010000010001101001110100001;
		#400 //-8.476653e-15 * -3.338003e-09 = 2.8295093e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100001101001001001011100101101;
		b = 32'b00011000111000101010000000011011;
		correct = 32'b10111011000100011011010001100110;
		#400 //-3.7951992e+20 * 5.8581296e-24 = -0.002223277
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000110100111111001101110100111;
		b = 32'b10110011100111101010110000010000;
		correct = 32'b10111010110001011101101010101111;
		#400 //20429.826 * -7.388746e-08 = -0.001509508
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011010011110001010000000010000;
		b = 32'b10101000111110010100110100010000;
		correct = 32'b10000011111100100001111010000111;
		#400 //5.1414495e-23 * -2.7677974e-14 = -1.423049e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111110000101101111000110111000;
		b = 32'b01000000001010010011100101101010;
		correct = 32'b01111110110001111000111011011010;
		#400 //5.015982e+37 * 2.6441293 = 1.3262905e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001100100010000010110101100011;
		b = 32'b11111110001000101001100110101100;
		correct = 32'b11001011001011001111110011101111;
		#400 //2.0981434e-31 * -5.403321e+37 = -11336943.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110100110100111011101000111101;
		b = 32'b10011011000001011110010111110010;
		correct = 32'b10010000010111010111101111011111;
		#400 //3.943732e-07 * -1.1075801e-22 = -4.3679992e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001111001100000111100110000110;
		b = 32'b10111110001111110011110010111101;
		correct = 32'b00001110000000111101010010001010;
		#400 //-8.7008745e-30 * -0.18675514 = 1.624933e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100011101101100000101001101111;
		b = 32'b11111101101101010100001000110000;
		correct = 32'b01100010000000001110010001110001;
		#400 //-1.9736898e-17 * -3.0116742e+37 = 5.9441104e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110010100001101001001100000000;
		b = 32'b10100010111111101011011100110001;
		correct = 32'b10010110000001011110011000100111;
		#400 //1.5666501e-08 * -6.90408e-18 = -1.0816278e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111111001111010101010110111110;
		b = 32'b10100111100111001100010101011001;
		correct = 32'b00100111011001111110010001101001;
		#400 //-0.7395896 * -4.3512663e-15 = 3.2181511e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101011110100010001110110111101;
		b = 32'b11001100011010100000111001011010;
		correct = 32'b01111000101111110011000011101000;
		#400 //-5.0561186e+26 * -61356390.0 = 3.102252e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001111000011101101101110100101;
		b = 32'b11111010010100000000011010111000;
		correct = 32'b11001001111010000010110001101100;
		#400 //7.0434425e-30 * -2.700335e+35 = -1901965.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011101110010000100001110100101;
		b = 32'b00111111001001001011111111011100;
		correct = 32'b00011101100000001110000101101100;
		#400 //5.30095e-21 * 0.64355254 = 3.41144e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101110011101110100101101100000;
		b = 32'b00101110001101011111010111100010;
		correct = 32'b00011101001011111100010111010000;
		#400 //5.6228244e-11 * 4.1373023e-11 = 2.3263324e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101111011101010010110110111100;
		b = 32'b01101000100100001011100100001000;
		correct = 32'b01011000100010101001101011101111;
		#400 //2.2298868e-10 * 5.467472e+24 = 1219184300000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111100011001110010100011101000;
		b = 32'b10000101010111010000110100011011;
		correct = 32'b01000010010001111001101000100110;
		#400 //-4.801001e+36 * -1.0393777e-35 = 49.900536
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101111100010100001100000001100;
		b = 32'b01001110101110101111111100010110;
		correct = 32'b01111110110010011011111000100101;
		#400 //8.5476e+28 * 1568639700.0 = 1.3408106e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010000100000010110010000110110;
		b = 32'b10111110001001001011000100000001;
		correct = 32'b10001111001001100111101101010011;
		#400 //5.103593e-29 * -0.16083147 = -8.208183e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100100111000001111101001000011;
		b = 32'b00100000100110111011010101010011;
		correct = 32'b01000110000010001101011011100000;
		#400 //3.3200831e+22 * 2.6378012e-19 = 8757.719
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110001011111100110000111011;
		b = 32'b00011000000101101101010111111011;
		correct = 32'b00010110110011110010100100111000;
		#400 //0.17167751 * 1.9495078e-24 = 3.3468666e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010011100000111100110001100101;
		b = 32'b01100001010101000011101001100000;
		correct = 32'b00110101010110101000011010100011;
		#400 //3.3270598e-27 * 2.4468226e+20 = 8.140725e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101001000110110011101110100110;
		b = 32'b00101011000111101110010001100110;
		correct = 32'b00010100110000001011001010011111;
		#400 //3.446865e-14 * 5.644984e-13 = 1.9457499e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000100000011000110010010111010;
		b = 32'b00010010000011101101001110100100;
		correct = 32'b10010110100111001010011111100000;
		#400 //-561.57385 * 4.5068167e-28 = -2.5309103e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100001101001101000100100101100;
		b = 32'b10111011010100011111011001110110;
		correct = 32'b00011101100010001001011001010001;
		#400 //-1.1284907e-18 * -0.0032037771 = 3.6154324e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101000100100111100101010010000;
		b = 32'b10100011111010110001111010011010;
		correct = 32'b11001101000001111011110010011101;
		#400 //5.583396e+24 * -2.5491711e-17 = -142330320.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111100111000101011101000001010;
		b = 32'b00111001101001100010010001100001;
		correct = 32'b00110111000100110010010011011011;
		#400 //0.027676601 * 0.00031689092 = 8.770464e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111011010000100001110110101010;
		b = 32'b00111110111000100000010111010110;
		correct = 32'b01111010101010110110001010011101;
		#400 //1.00790725e+36 * 0.44145077 = 4.4494144e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111110010000011011101110111110;
		b = 32'b01110101000111101010110011001100;
		correct = 32'b11110011111100000010100101001000;
		#400 //-0.18919274 * 2.0114444e+32 = -3.805507e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100000110100010010011011111011;
		b = 32'b01111100100101011000011001101001;
		correct = 32'b11011101111101000101001100000001;
		#400 //-3.5431772e-19 * 6.211027e+36 = -2.200677e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110011000110110000110101110100;
		b = 32'b01000010011010111010001110010100;
		correct = 32'b10110110000011101011100001101101;
		#400 //-3.6100985e-08 * 58.909744 = -2.1266999e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101100110100011000001010000001;
		b = 32'b10110011100110111110100101111000;
		correct = 32'b11100000111111110011001000101100;
		#400 //2.0262543e+27 * -7.260218e-08 = -1.4711047e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011110111111111110010110111000;
		b = 32'b00100000100101000111010001110000;
		correct = 32'b11000000000101000110010100110010;
		#400 //-9.2196733e+18 * 2.5149227e-19 = -2.3186765
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010101111010111000100001010111;
		b = 32'b11011000010101101100111011110000;
		correct = 32'b11101110110001011010001001011101;
		#400 //32371350000000.0 * -944737100000000.0 = -3.0582416e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100101000111011111100101011011;
		b = 32'b01001110010110011101011001000111;
		correct = 32'b10110100000001100110110010011000;
		#400 //-1.3702064e-16 * 913674700.0 = -1.2519229e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011110011111111100100100010111;
		b = 32'b00000011101111011010010001010000;
		correct = 32'b10100010101111010111101110100011;
		#400 //-4.607822e+18 * 1.1146146e-36 = -5.135946e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001100111110001111111011001111;
		b = 32'b00100111110101110011000100111110;
		correct = 32'b00110101010100010100110111100101;
		#400 //130545270.0 * 5.9727876e-15 = 7.797192e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001100100100001011011011011100;
		b = 32'b00111001011100111000010010111001;
		correct = 32'b10000110100010011010100010011010;
		#400 //-2.2296767e-31 * 0.00023223729 = -5.178141e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001010001100101011001010100011;
		b = 32'b00111000001011100101111110010110;
		correct = 32'b00000010111100110111000001001000;
		#400 //8.603986e-33 * 4.1573854e-05 = 3.5770087e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100110000101101110101100000100;
		b = 32'b00110000010000111110101110110000;
		correct = 32'b10010110111001101111111111101011;
		#400 //-5.236021e-16 * 7.127552e-10 = -3.732001e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011100100011011111111101001010;
		b = 32'b01100000000011010100101000001010;
		correct = 32'b00111101000111001011110101011010;
		#400 //9.396588e-22 * 4.0723844e+19 = 0.038266517
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001100010000011101001001101111;
		b = 32'b11110011011100111010100000000001;
		correct = 32'b11000000001110000111100111110010;
		#400 //1.4931504e-31 * -1.9304438e+31 = -2.882443
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011110100011111101011001000011;
		b = 32'b11000011001000111000000100001110;
		correct = 32'b11100010001101111011101111011111;
		#400 //5.1822726e+18 * -163.50412 = -8.473229e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111000100110111011010110101110;
		b = 32'b01101101000100110010110010111011;
		correct = 32'b11100110001100110000100100010000;
		#400 //-7.4248164e-05 * 2.8467733e+27 = -2.113677e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110010011110101101101001000100;
		b = 32'b01001001110001111000111001000101;
		correct = 32'b10111100110000111000101100010100;
		#400 //-1.4601543e-08 * 1634760.6 = -0.023870029
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000000001001000110110111110011;
		b = 32'b00100101001011010111001010011010;
		correct = 32'b00100101110111101100111111010010;
		#400 //2.5692108 * 1.5044187e-16 = 3.8651686e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110011110100111100110101000110;
		b = 32'b10010111001101101000001101110110;
		correct = 32'b00001011100101110000000010110011;
		#400 //-9.862792e-08 * -5.89733e-25 = 5.8164136e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100000101000101000100100110111;
		b = 32'b11001101011010001000110010010101;
		correct = 32'b01101110100100111010010110011011;
		#400 //-9.369562e+19 * -243845460.0 = 2.284725e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111011100010001000111100001000;
		b = 32'b10101011101010101001001111010111;
		correct = 32'b11100111101101011111101110110000;
		#400 //1.4181068e+36 * -1.212026e-12 = -1.7187823e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010101100110111010011100101100;
		b = 32'b10110101000101111000101001000000;
		correct = 32'b00001011001110000100011101010100;
		#400 //-6.286775e-26 * -5.6453064e-07 = 3.5490772e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000011011110101101011010100110;
		b = 32'b01001110100011110010101010100111;
		correct = 32'b00010010100011000100011110110010;
		#400 //7.37148e-37 * 1200968600.0 = 8.852916e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110011011000001000000010011001;
		b = 32'b01101000101111100000000101011001;
		correct = 32'b01011100101001101010000010100000;
		#400 //5.2271023e-08 * 7.178196e+24 = 3.7521164e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110101100100100100010010110001;
		b = 32'b01110000101010010110101011111110;
		correct = 32'b11100110110000011001100011110101;
		#400 //-1.089784e-06 * 4.194585e+29 = -4.5711915e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110111000101000100010011000;
		b = 32'b00110110010111110101111110010000;
		correct = 32'b10101101110001011010100110001101;
		#400 //-6.7512265e-06 * 3.3285214e-06 = -2.2471603e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110101110011001100010100111010;
		b = 32'b00100000111011110000001011000110;
		correct = 32'b11010111001111110010111001011001;
		#400 //-5.191547e+32 * 4.049001e-19 = -210205780000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100011110011101011110101100001;
		b = 32'b10001010101000111110001111010110;
		correct = 32'b10101111000001000101101010010100;
		#400 //7.627351e+21 * -1.5782031e-32 = -1.203751e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100100000101001001101010010100;
		b = 32'b10101010111011000100010001011010;
		correct = 32'b10001111100010010010011000101110;
		#400 //3.2223317e-17 * -4.196945e-13 = -1.352395e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001110001001100110101111010000;
		b = 32'b00011001110110010010001110101111;
		correct = 32'b10101000100011010010100010010110;
		#400 //-698020860.0 * 2.2451687e-23 = -1.5671746e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011001010011101101011010111000;
		b = 32'b00101110010111011110000111101101;
		correct = 32'b11001000001100110100010111100111;
		#400 //-3638745700000000.0 * 5.0450245e-11 = -183575.61
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000011000101011111101101000111;
		b = 32'b00111110000000010100011000110101;
		correct = 32'b00000001100101110111100110000001;
		#400 //4.4075617e-37 * 0.12624438 = 5.564299e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001010011011111010111100001110;
		b = 32'b10100101101110011010110100010001;
		correct = 32'b00110000101011011101011110001010;
		#400 //-3926979.5 * -3.2209659e-16 = 1.2648667e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001111011100011001011010111110;
		b = 32'b11001111010011111011010111000110;
		correct = 32'b01011111010001000000010001101110;
		#400 //-4053188000.0 * -3484796400.0 = 1.4124535e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100111011100111101010111010101;
		b = 32'b01111000101001100001100001100010;
		correct = 32'b01100000100111100011001111100010;
		#400 //3.3838943e-15 * 2.6950494e+34 = 9.119763e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111111100011111001000111000101;
		b = 32'b10001100001000110100011011111101;
		correct = 32'b10001100001101110010001101000000;
		#400 //1.121636 * -1.2578425e-31 = -1.4108415e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010000011111111110011011011010;
		b = 32'b01101100000100110001011111110000;
		correct = 32'b00111101000100110000100101111101;
		#400 //5.0467724e-29 * 7.1130055e+26 = 0.03589772
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011101111010100011000100000010;
		b = 32'b10011111100010101101111110001110;
		correct = 32'b10111101111111100001010111011011;
		#400 //2.109409e+18 * -5.8815114e-20 = -0.12406512
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011100011101101101001010010001;
		b = 32'b00010000001000011001000100101111;
		correct = 32'b00101101000110111100011001101000;
		#400 //2.7789746e+17 * 3.1863497e-29 = 8.854785e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000101000011010110101011111100;
		b = 32'b10011010000010111101111010011000;
		correct = 32'b00011111100110101000100000011011;
		#400 //-2262.6865 * -2.8924336e-23 = 6.5446705e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110110000111110111011000101011;
		b = 32'b00000100110001011010010001100110;
		correct = 32'b10111011011101100011100010101101;
		#400 //-8.0856634e+32 * 4.6465454e-36 = -0.0037570402
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101111001111110010111101000010;
		b = 32'b00011010010100010100011111111010;
		correct = 32'b01001010000111000100101101010110;
		#400 //5.916877e+28 * 4.327833e-23 = 2560725.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111000001111010110111011001100;
		b = 32'b01000001100111111101001101101111;
		correct = 32'b01111010011011001000100010001010;
		#400 //1.5368615e+34 * 19.97824 = 3.0703785e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011101000101111111100100011111;
		b = 32'b01001101101100011111110110000011;
		correct = 32'b00101011010100110101001101111011;
		#400 //2.0113476e-21 * 373272670.0 = 7.507811e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111000010100010011001110110110;
		b = 32'b10101001001101111010011011101001;
		correct = 32'b11100010000101100001010001011101;
		#400 //1.6972482e+34 * -4.0778934e-14 = -6.921197e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011111111101110011000011101111;
		b = 32'b10100110111101011010001001000011;
		correct = 32'b10000111011011010010111010000010;
		#400 //1.0468952e-19 * -1.7044271e-15 = -1.7843566e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100000010101111011010011101110;
		b = 32'b01010000110101101110101100111000;
		correct = 32'b11110001101101010001011101110001;
		#400 //-6.217324e+19 * 28845916000.0 = -1.793444e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101010100001000101011110101101;
		b = 32'b01010011001010001011110001010011;
		correct = 32'b11111110001011100111010111001010;
		#400 //-7.999612e+25 * 724714060000.0 = -5.7974317e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011110010111101011110110000000;
		b = 32'b11000110011010010100011111011011;
		correct = 32'b01100101010010101111100011111111;
		#400 //-4.0125313e+18 * -14929.964 = 5.990695e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111010001011100000000010110001;
		b = 32'b10001001101101100111001110011110;
		correct = 32'b10000100011110000000011000100111;
		#400 //0.0006637676 * -4.3923632e-33 = -2.9155085e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111001100110100010100000011000;
		b = 32'b00100000110010001110011011000110;
		correct = 32'b10011010111100011111010010010100;
		#400 //-0.0002940304 * 3.403403e-19 = -1.000704e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111111111101110000110101100101;
		b = 32'b11101001011001101111101100100001;
		correct = 32'b11111111111101110000110101100101;
		#400 //nan * -1.7452429e+25 = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110110001011010010111001110010;
		b = 32'b11100110000111001100111011011011;
		correct = 32'b11011100110101000010100001111010;
		#400 //2.5806044e-06 * -1.8512625e+23 = -4.777376e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010110101100011011101011110111;
		b = 32'b01100000111001001101000001001100;
		correct = 32'b01111000000111101101101100100001;
		#400 //97708280000000.0 * 1.3190209e+20 = 1.2887928e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001010011010111011000111001011;
		b = 32'b01001000001111101100110000001110;
		correct = 32'b01010011001011111010100111010011;
		#400 //3861618.8 * 195376.22 = 754468450000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000111000001011111100111110001;
		b = 32'b10110010010111011001000101010010;
		correct = 32'b00111001111001111110100110100101;
		#400 //-34297.94 * -1.2896935e-08 = 0.00044233832
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100000101111111000110111101010;
		b = 32'b10110000101100011010110111100010;
		correct = 32'b00010010000001001111001100111011;
		#400 //-3.245057e-19 * -1.2927865e-09 = 4.195166e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111011111001110111000101101101;
		b = 32'b00011011111001110110110000010001;
		correct = 32'b10011000010100010011100100001101;
		#400 //-0.007063082 * 3.828558e-22 = -2.704142e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100111110100101010001010011111;
		b = 32'b00110110101101010111100001110110;
		correct = 32'b10011111000101010101000000011000;
		#400 //-5.8463023e-15 * 5.408244e-06 = -3.161823e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011100000100110111011011001111;
		b = 32'b00001110001010101100000011110000;
		correct = 32'b00101010110001001011100000010010;
		#400 //1.6602981e+17 * 2.1047014e-30 = 3.4944318e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111000010100101010011110101001;
		b = 32'b00011000000101110000000101101100;
		correct = 32'b10010000111110001000010000100000;
		#400 //-5.0224047e-05 * 1.951701e-24 = -9.8022323e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100000111001001000010110010011;
		b = 32'b00001111010001011110110000101100;
		correct = 32'b10110000101100001010110110011101;
		#400 //-1.3173383e+20 * 9.758335e-30 = -1.2855029e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110000000011100100011001110;
		b = 32'b00001001000110001000110011011011;
		correct = 32'b00000111100110101010110101000110;
		#400 //0.12674257 * 1.8362564e-33 = 2.3273186e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100110111010100100011110010100;
		b = 32'b11000111101011101011111001110000;
		correct = 32'b00101111000111111110101011101110;
		#400 //-1.6256413e-15 * -89468.875 = 1.454443e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110110010111100110111101010001;
		b = 32'b00011001101101110001111110100100;
		correct = 32'b01010000100111110001110100010001;
		#400 //1.1278786e+33 * 1.8934536e-23 = 21355858000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100000011111001001011111100100;
		b = 32'b10011101100001101001111001111000;
		correct = 32'b00111110100001001101001111011101;
		#400 //-7.280507e+19 * -3.5633358e-21 = 0.2594289
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011011101000110000001011110111;
		b = 32'b11110000001001001011011001110110;
		correct = 32'b01001100010100011100010000101011;
		#400 //-2.6968004e-22 * -2.039045e+29 = 54988972.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001111100110100010010100011010;
		b = 32'b10111001111100010100011111011110;
		correct = 32'b11001010000100010100100000110011;
		#400 //5172245500.0 * -0.00046020647 = -2380300.8
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100001111010000100111001111000;
		b = 32'b00000101010011110000100001001111;
		correct = 32'b00100111101110111101111011111101;
		#400 //5.3566236e+20 * 9.734619e-36 = 5.214469e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100111011001010111001111111101;
		b = 32'b10110010001000001100100010111101;
		correct = 32'b11011010000100000001110001101010;
		#400 //1.0835615e+24 * -9.358868e-09 = -1.014091e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010011001001111100110001010110;
		b = 32'b01100000101001000000110100111110;
		correct = 32'b11110100010101110000111100101010;
		#400 //-720687700000.0 * 9.456938e+19 = -6.815499e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000001000101001011110110010101;
		b = 32'b01100001110010001101101010110101;
		correct = 32'b10100011011010010110011001011110;
		#400 //-2.7319325e-38 * 4.6313854e+20 = -1.2652632e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100101010000000101110000010110;
		b = 32'b11111000100110111100011001101001;
		correct = 32'b11011110011010100001100110101111;
		#400 //1.6684545e-16 * -2.5275945e+34 = -4.2171766e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000010000000010110000000110011;
		b = 32'b00010000101101011101101100011011;
		correct = 32'b00010011001101111100111101111110;
		#400 //32.343945 * 7.17295e-29 = 2.3200149e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111101100100110101101001011100;
		b = 32'b00011110111110100100010111000000;
		correct = 32'b11011101000100000000111001100100;
		#400 //-2.448321e+37 * 2.6498628e-20 = -6.487715e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101100100101101100001110010101;
		b = 32'b11101110010011101011001101011101;
		correct = 32'b11011011011100110111011000000111;
		#400 //4.2849704e-12 * -1.5992687e+28 = -6.852819e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011010101010011100100011000110;
		b = 32'b11110111101110110111101101000111;
		correct = 32'b11010010111110001010111011010110;
		#400 //7.022113e-23 * -7.605155e+33 = -534042570000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110100010010101100110011101101;
		b = 32'b10111111011001110011011001000010;
		correct = 32'b11110100001101110010100111100101;
		#400 //6.427004e+31 * -0.90317166 = -5.804688e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100000111101000110110011001011;
		b = 32'b01001111110100100101010111101100;
		correct = 32'b00110001010010001101001101001000;
		#400 //4.14072e-19 * 7057692700.0 = 2.922393e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011011011100100101010011100011;
		b = 32'b00001110101101000111010111100111;
		correct = 32'b10101010101010101101001101001011;
		#400 //-6.821028e+16 * 4.448696e-30 = -3.034468e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111111000011101100000010110010;
		b = 32'b00001101010111011010011101001010;
		correct = 32'b01001100111101110011001101000101;
		#400 //1.897509e+38 * 6.830225e-31 = 129604136.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110000011111111101011111000101;
		b = 32'b00100011100110111111111111010001;
		correct = 32'b01010100100110111110011101001101;
		#400 //3.167181e+29 * 1.6913476e-17 = 5356804000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001000011110011011101010001001;
		b = 32'b10010010010000011111110111101110;
		correct = 32'b00011011001111010011110101010111;
		#400 //-255722.14 * -6.1213054e-28 = 1.5653534e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011011001000011011001001100110;
		b = 32'b11101000000110111011000001101011;
		correct = 32'b11000011110001001010110011100100;
		#400 //1.3375252e-22 * -2.9408846e+24 = -393.3507
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100100111010100011111111010;
		b = 32'b00100001001010100110000011101011;
		correct = 32'b00100110010100010101101010101111;
		#400 //1258.2493 * 5.772651e-19 = 7.263434e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111011110110000101101011000001;
		b = 32'b00010001010000000001000000000101;
		correct = 32'b00001101101000100101000110011011;
		#400 //0.0066026156 * 1.5151066e-28 = 1.0003667e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011111110110111000101100101101;
		b = 32'b00111101000001111000011001100011;
		correct = 32'b10011101011010000111001101001001;
		#400 //-9.2980355e-20 * 0.033087146 = -3.0764545e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010110111011110000111110000100;
		b = 32'b01000111001001110100111100101000;
		correct = 32'b01011110100111000011110100001010;
		#400 //131424960000000.0 * 42831.156 = 5.629083e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010011111001110111000011111101;
		b = 32'b01101001100011001100100001101010;
		correct = 32'b01111101111111101000110111110101;
		#400 //1988066100000.0 * 2.1274505e+25 = 4.2295124e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000001111000011110110000111000;
		b = 32'b00101110011000010001010111011101;
		correct = 32'b00110000110001101010001111101001;
		#400 //28.240341 * 5.1178495e-11 = 1.4452982e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101100001010100001111101110000;
		b = 32'b00110110100100011000110100101001;
		correct = 32'b01100011010000010111001100111010;
		#400 //8.226634e+26 * 4.33777e-06 = 3.5685246e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111011010001010010000101000110;
		b = 32'b01010100110111100101001011000110;
		correct = 32'b11010000101010110011001010011000;
		#400 //-0.0030079647 * 7638971600000.0 = -22977757000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001100100111011000111110001011;
		b = 32'b11010100110001010010111011011111;
		correct = 32'b00100001111100101011100010011110;
		#400 //-2.4276072e-31 * -6775159400000.0 = 1.6447426e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011101111111001111011101001100;
		b = 32'b01000010000101000010101110010001;
		correct = 32'b00100000100100100110101000000101;
		#400 //6.6959544e-21 * 37.042545 = 2.480352e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010100001101011010101011000111;
		b = 32'b01101110000100101011001011101010;
		correct = 32'b01000010110100000011010010111001;
		#400 //9.171845e-27 * 1.1350276e+28 = 104.102974
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000101111001101101011111110100;
		b = 32'b11101010100011111101011010101100;
		correct = 32'b10110001000000011011010000110101;
		#400 //2.1708425e-35 * -8.694508e+25 = -1.8874406e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011000101011000110101110000001;
		b = 32'b11001110010100100000110111110101;
		correct = 32'b11100111100011010111100110010110;
		#400 //1516621800000000.0 * -881032500.0 = -1.3361931e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010101100010101111111001011110;
		b = 32'b11100101101011011001001000001101;
		correct = 32'b00111011101111000111101001100011;
		#400 //-5.6139077e-26 * -1.02457945e+23 = 0.0057518943
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111110100011001010010100010001;
		b = 32'b00001011000000010011011110111011;
		correct = 32'b11001010000011011111101110011000;
		#400 //-9.34745e+37 * 2.4886423e-32 = -2326246.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010110110111000110111001000011;
		b = 32'b00101011010100010100011110101001;
		correct = 32'b01000010101101000011001110111001;
		#400 //121183064000000.0 * 7.4351164e-13 = 90.10102
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100111100101010010010110010101;
		b = 32'b00100101100100110011010111111110;
		correct = 32'b11001101101010111000100000010011;
		#400 //-1.4086517e+24 * 2.5537022e-16 = -359727700.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100011001111100010100101111111;
		b = 32'b11110100110010100111010000110010;
		correct = 32'b11011000100101100110001100001110;
		#400 //1.0308708e-17 * -1.283204e+32 = -1322817400000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110010000010111001100111101101;
		b = 32'b00010111110101110010000011101010;
		correct = 32'b00001010011010101010000001110010;
		#400 //8.1258635e-09 * 1.3902358e-24 = 1.12968666e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100010110001001101001010001100;
		b = 32'b01010011101010110001110111101110;
		correct = 32'b10110111000000111000111110100110;
		#400 //-5.334883e-18 * 1469883100000.0 = -7.841654e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001101010011110001001010100101;
		b = 32'b11010001000101101011101101110100;
		correct = 32'b10011110111100111101100100011010;
		#400 //6.380924e-31 * -40461877000.0 = -2.5818417e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011110110111101100000100110101;
		b = 32'b10111011001110010010001011011000;
		correct = 32'b11011010101000010001011111110001;
		#400 //8.0255844e+18 * -0.0028249528 = -2.2671898e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101011110000100000111001101101;
		b = 32'b11010101100111100001010000001010;
		correct = 32'b01000001111011111010100000110000;
		#400 //-1.3788533e-12 * -21726113000000.0 = 29.957123
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001000101001101100110111101011;
		b = 32'b01111101011000110000001110101001;
		correct = 32'b01000110100100111110101011111010;
		#400 //1.0039173e-33 * 1.885961e+37 = 18933.488
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011110010110101010111000111110;
		b = 32'b01011001001101000011011101101001;
		correct = 32'b00111000000110011111000111011001;
		#400 //1.1576856e-20 * 3170401200000000.0 = 3.670328e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111011000011101110110001110001;
		b = 32'b11110011011010111001110010101000;
		correct = 32'b01101111000000111000101010000010;
		#400 //-0.002180841 * -1.8667101e+31 = 4.070998e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001111001010001000100101110001;
		b = 32'b11000010111110110100010011011100;
		correct = 32'b11010010101001010110110000010111;
		#400 //2827579600.0 * -125.63449 = -355241530000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110101000111111001111111100001;
		b = 32'b11111101011110101001111101111110;
		correct = 32'b11110011000111000100010110010101;
		#400 //5.946477e-07 * -2.0820946e+37 = -1.2381128e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000000110010000010100111111011;
		b = 32'b10111111100100011101011000100001;
		correct = 32'b11000000111001000000111001101000;
		#400 //6.2551246 * -1.1393472 = -7.1267586
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110101101110111101100101011011;
		b = 32'b01101100111011101111100101011111;
		correct = 32'b11100011001011110101101100001111;
		#400 //-1.3995844e-06 * 2.3112157e+27 = -3.2347417e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000010010010001100100000001000;
		b = 32'b10101011110100101111111000001111;
		correct = 32'b10101110101001010111101101011001;
		#400 //50.195343 * -1.4991913e-12 = -7.525242e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101001101111111001100110011111;
		b = 32'b00111101100101100001111100001000;
		correct = 32'b00100111111000001011011001111010;
		#400 //8.508753e-14 * 0.073301375 = 6.237033e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001100011110110011011011001110;
		b = 32'b10111111001100010011100011010000;
		correct = 32'b00001100001011011110100010100101;
		#400 //-1.9352829e-31 * -0.69227314 = 1.3397444e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010100111110111111100101100111;
		b = 32'b00110100010000101111100011101110;
		correct = 32'b00001001101111111110100000000100;
		#400 //2.5442895e-26 * 1.8158218e-07 = 4.6199764e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001100100010111010101101000010;
		b = 32'b10010010010000100000110111110011;
		correct = 32'b10011111010100111011111011001001;
		#400 //73226770.0 * -6.12328e-28 = -4.4838802e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010001101111110011010011111011;
		b = 32'b00111111010111100000110111011010;
		correct = 32'b10010001101001011101101001001010;
		#400 //-3.0167138e-28 * 0.86739886 = -2.616694e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110011001110110101010011101001;
		b = 32'b11110111010001110001010000011011;
		correct = 32'b11101011000100011010110110111000;
		#400 //4.3616556e-08 * -4.0377924e+33 = -1.761146e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001000101100001000001111111101;
		b = 32'b11001001111101001000000000011100;
		correct = 32'b00010011001010001001011000100010;
		#400 //-1.0623645e-33 * -2002947.5 = 2.1278602e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101110101011010101110011011000;
		b = 32'b00111101011001000111110001111100;
		correct = 32'b11101100100110101011101011111101;
		#400 //-2.6826574e+28 * 0.05578278 = -1.4964608e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010001001010001111100100000001;
		b = 32'b10000100110001101000111000011111;
		correct = 32'b00010110100000110000111001100101;
		#400 //-45358256000.0 * -4.6680094e-36 = 2.1173276e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100101101111100000010101001001;
		b = 32'b11010010100101000000110011111010;
		correct = 32'b10111000110110111100100101100000;
		#400 //3.2963327e-16 * -317936440000.0 = -0.00010480243
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000000111011010101011001110000;
		b = 32'b01000101100010111001010100101001;
		correct = 32'b11000111000000010110100000111000;
		#400 //-7.4168015 * 4466.645 = -33128.22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101010010000111111100000010011;
		b = 32'b01110111011000011110010000101110;
		correct = 32'b11100010001011001110101110110101;
		#400 //-1.7405547e-13 * 4.5816204e+33 = -7.974561e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100111110101101010100010101010;
		b = 32'b01000100110001110111110010011100;
		correct = 32'b01101101001001110100010110011001;
		#400 //2.0273955e+24 * 1595.894 = 3.2355084e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101001100110111011000101010010;
		b = 32'b10011011100111010010000001000000;
		correct = 32'b10000101101111110001111010111001;
		#400 //6.914143e-14 * -2.5994312e-22 = -1.797284e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000110000011010111100010110000;
		b = 32'b00000001111001011010001010001010;
		correct = 32'b00001000011111011100110110010000;
		#400 //9054.172 * 8.4354547e-38 = 7.6376056e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011111011001101011000001101010;
		b = 32'b00100001110001101000101100000010;
		correct = 32'b01000001101100101110100110110110;
		#400 //1.6622903e+19 * 1.3453797e-18 = 22.364117
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101101100110000011100001101110;
		b = 32'b00111000101100010001011101010101;
		correct = 32'b00100110110100101001100111000111;
		#400 //1.730546e-11 * 8.4443636e-05 = 1.4613359e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100110010000111111111101100011;
		b = 32'b10001100110110010011000101010011;
		correct = 32'b00110011101001100100100100111110;
		#400 //-2.3139313e+23 * -3.346383e-31 = 7.7433e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101101010100011010000010101000;
		b = 32'b10011101001000101010001111111110;
		correct = 32'b00001011000001010010110111110100;
		#400 //-1.1915947e-11 * -2.1525303e-21 = 2.564944e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100010100000101110000000001;
		b = 32'b11100011001111110000101100100110;
		correct = 32'b11101000000110110111110110111000;
		#400 //833.43756 * -3.5241314e+21 = -2.9371436e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010110000011000100001101110110;
		b = 32'b00111101100110111101010101101001;
		correct = 32'b00010100001010101100001110001100;
		#400 //1.1330397e-25 * 0.07609064 = 8.6213715e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100101000110110111011111000101;
		b = 32'b01001111111000100000101101100011;
		correct = 32'b01110101100010010100011010100110;
		#400 //4.588601e+22 * 7584794000.0 = 3.4803593e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101110110010101001110111000111;
		b = 32'b00001100010110101100010110000110;
		correct = 32'b00111011101011010010011010110001;
		#400 //3.1353357e+28 * 1.6853549e-31 = 0.0052841534
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100110001010010011011011100000;
		b = 32'b11100001101001100101101101011101;
		correct = 32'b01001000010110111110101111110010;
		#400 //-5.8708023e-16 * -3.8359287e+20 = 225199.78
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010001111100011100000011000000;
		b = 32'b01101001011101000111101100001110;
		correct = 32'b00111011111001101101111111101100;
		#400 //3.8141887e-28 * 1.8472438e+25 = 0.0070457365
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100100010100000001110000111000;
		b = 32'b11011100110011000100111010110010;
		correct = 32'b11000001101001100001011001110110;
		#400 //4.5126713e-17 * -4.6005937e+17 = -20.760967
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000110100011010111001001000110;
		b = 32'b00001001110011101100000100111110;
		correct = 32'b10010000111001000111100101110011;
		#400 //-18105.137 * 4.977442e-33 = -9.0117265e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111001001111000011000001101010;
		b = 32'b10010100100011100100110100111110;
		correct = 32'b11001110010100010011011101000110;
		#400 //6.107086e+34 * -1.4368802e-26 = -877515140.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011000110001100001011100111010;
		b = 32'b11000111101010101111111101101011;
		correct = 32'b11100001000001000101000100010000;
		#400 //1742424500000000.0 * -87550.836 = -1.5255071e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011000000000101001000111000100;
		b = 32'b01111101100110110111010110000110;
		correct = 32'b11010110000111101001010001100101;
		#400 //-1.68757e-24 * 2.583007e+37 = -43590047000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111000001110110001110110010111;
		b = 32'b10100011001001101110110010110101;
		correct = 32'b10011011111101000000010001100111;
		#400 //4.4611832e-05 * -9.049003e-18 = -4.036926e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101011110111111100110000010100;
		b = 32'b00111010001000111110001110010000;
		correct = 32'b01100110100011110100010111100001;
		#400 //5.4110838e+26 * 0.0006251866 = 3.3829372e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111100110001101001000100011100;
		b = 32'b10001100010111110110011100101011;
		correct = 32'b01001001101011010100100001101101;
		#400 //-8.2481436e+36 * -1.7210341e-31 = 1419533.6
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110000111000100010010000011000;
		b = 32'b10101001011100010101010011110111;
		correct = 32'b01011010110101010010111100001001;
		#400 //-5.5989798e+29 * -5.3586445e-14 = 3.0002943e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010011000110010011000011110011;
		b = 32'b10110010110000101111111100011100;
		correct = 32'b11000110011010010101111110000001;
		#400 //657951200000.0 * -2.2700583e-08 = -14935.876
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011101100101101000011100000000;
		b = 32'b11010110101010110101001100111111;
		correct = 32'b11110100110010010111101001000000;
		#400 //1.3558298e+18 * -94187010000000.0 = -1.2770156e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001001101001101110001001101001;
		b = 32'b01001101110010111001001111101001;
		correct = 32'b11011000000001001011010111110101;
		#400 //-1367117.1 * 426933540.0 = -583668140000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101011101101010011010100000010;
		b = 32'b00000011011101110100010011101000;
		correct = 32'b10101111101011110000011011101011;
		#400 //-4.381318e+26 * 7.2665877e-37 = -3.183723e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001110001010011011111010001010;
		b = 32'b11101111111000000010001000111001;
		correct = 32'b11111110100101001001110101101010;
		#400 //711959200.0 * -1.3873203e+29 = -9.877154e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100010100111000010011001001101;
		b = 32'b10110010001111111010100000001011;
		correct = 32'b00010101011010011100111000100111;
		#400 //-4.2324437e-18 * -1.1155872e-08 = 4.72166e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010110011100001110110011111001;
		b = 32'b00100011001010010101001011011111;
		correct = 32'b10111010000111110101101001101110;
		#400 //-66225145000000.0 * 9.179057e-18 = -0.0006078844
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110001000101001011111010001110;
		b = 32'b11101101000100101011111001100100;
		correct = 32'b01011110101010101000011010011001;
		#400 //-2.1645152e-09 * -2.8384362e+27 = 6.1438384e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111011001101111000101101010100;
		b = 32'b10001100100000100000111111101010;
		correct = 32'b11001000001110101000000001010011;
		#400 //9.530162e+35 * -2.003925e-31 = -190977.3
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110100100100111110001101101100;
		b = 32'b10111111011110010101100100001110;
		correct = 32'b10110100100100000000101110100110;
		#400 //2.7546355e-07 * -0.9740151 = -2.6830566e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110000000000100100001010010010;
		b = 32'b00010010110110000010100001100101;
		correct = 32'b00000011010110111111100101110010;
		#400 //4.7388327e-10 * 1.3641474e-27 = 6.4644665e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110010011001010100001001011010;
		b = 32'b10011101100100001111100100111111;
		correct = 32'b11010000100000011101010010001001;
		#400 //4.540946e+30 * -3.8374197e-21 = -17425517000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101010110101001011111001110010;
		b = 32'b11100101001101011001011010111000;
		correct = 32'b11010000100101101110011111100111;
		#400 //3.7790913e-13 * -5.3595538e+22 = -20254243000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100010110111110111111010110000;
		b = 32'b10110100101110111101010000000011;
		correct = 32'b00011000001000111111101010100010;
		#400 //-6.0578407e-18 * -3.4985723e-07 = 2.1193793e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110011000101111101110111100;
		b = 32'b10100000010101001001011100011000;
		correct = 32'b00010111001111000111111001101111;
		#400 //-3.3823153e-06 * -1.8007091e-19 = 6.090566e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101011101101100110101101000110;
		b = 32'b10111000011001101111011001110011;
		correct = 32'b01100100101001001001001111111110;
		#400 //-4.4106217e+26 * -5.5065797e-05 = 2.428744e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011001010001001010010000010010;
		b = 32'b11001111100010010111110010101001;
		correct = 32'b01101001010100110011011100011110;
		#400 //-3459343300000000.0 * -4613296600.0 = 1.5958977e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011100001110110101111111011011;
		b = 32'b11000111001100001101101100011000;
		correct = 32'b10100100000000010111001001000011;
		#400 //6.1997e-22 * -45275.094 = -2.80692e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101101110111001101110000100100;
		b = 32'b01000010001011001010111100000001;
		correct = 32'b10110000100101001111101011100100;
		#400 //-2.5108866e-11 * 43.170902 = -1.0839725e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110101100110001101000110011101;
		b = 32'b00010100010000001000010000110001;
		correct = 32'b11001010011001011101100000111110;
		#400 //-3.874417e+32 * 9.719593e-27 = -3765775.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011110000110100001111000011100;
		b = 32'b10000100100100100001010011100000;
		correct = 32'b10100011001011111110001101111010;
		#400 //2.776336e+18 * -3.4343606e-36 = -9.534939e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101000011010011011101110111000;
		b = 32'b10000111110111000101011000110001;
		correct = 32'b00110000110010010010110000000100;
		#400 //-4.4150968e+24 * -3.315258e-34 = 1.4637185e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000000111111111000000011001100;
		b = 32'b11000110001101010110110001100110;
		correct = 32'b01000111101101010001001001000000;
		#400 //-7.9844723 * -11611.1 = 92708.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010111010001000110011011010001;
		b = 32'b00001111101110110011001011001110;
		correct = 32'b00100111100011111001111000010101;
		#400 //215945870000000.0 * 1.8459193e-29 = 3.9861866e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110100111010110110000111100100;
		b = 32'b00110111110101100101010111000001;
		correct = 32'b00101101010001010001001010101110;
		#400 //4.3843386e-07 * 2.555072e-05 = 1.1202301e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011001001011000101100011000010;
		b = 32'b00111111001000110100111101011010;
		correct = 32'b01011000110110111110001111011111;
		#400 //3031955400000000.0 * 0.63792956 = 1934174000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011011011101010101110010001110;
		b = 32'b00110011111111001000101001000110;
		correct = 32'b11001111111100100000101110100011;
		#400 //-6.9063134e+16 * 1.1759816e-07 = -8121698000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111001000010011111100001111101;
		b = 32'b10111100110111111011101001001001;
		correct = 32'b01110110011100010010011110110110;
		#400 //-4.477404e+34 * -0.027310507 = 1.2228017e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000001001110101010101100111110;
		b = 32'b01110001000000000101011101100100;
		correct = 32'b11110010101110110010101010110000;
		#400 //-11.666807 * 6.355157e+29 = -7.414439e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001110100001001000100001100000;
		b = 32'b11000000101001110111111011000111;
		correct = 32'b01001111101011010110110100110010;
		#400 //-1111765000.0 * -5.2342257 = 5819229000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001100000101101111001100111101;
		b = 32'b01100001111110100110111100101011;
		correct = 32'b10101110100100111010101100010110;
		#400 //-1.1628777e-31 * 5.7746206e+20 = -6.715177e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111111010111100110100100010001;
		b = 32'b00101110100000101111011000000100;
		correct = 32'b10101110011000111000111000101110;
		#400 //-0.8687907 * 5.955417e-11 = -5.1740105e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100101011100010000011000000000;
		b = 32'b10110000101010000111010100101001;
		correct = 32'b11010110100111101001101000111110;
		#400 //7.1137563e+22 * -1.2256908e-09 = -87192650000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100000110000010010100100100000;
		b = 32'b10011001000100011100001101000101;
		correct = 32'b00111010010110111111011101000011;
		#400 //-1.1134953e+20 * -7.535759e-24 = 0.0008391032
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000001000011111110000010110100;
		b = 32'b01011011110101101111001001001010;
		correct = 32'b01011101011100011001110000000101;
		#400 //8.992359 * 1.2100409e+17 = 1.08811223e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010010101010011011111111101110;
		b = 32'b10111011011000100011010000100100;
		correct = 32'b11001110100101011111111000000011;
		#400 //364534760000.0 * -0.0034515942 = -1258226000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010000100000101010000101110001;
		b = 32'b11011000001010011001010100110110;
		correct = 32'b10101001001011010001000101101110;
		#400 //5.15247e-29 * -745833300000000.0 = -3.8428834e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000101100001110101110011101101;
		b = 32'b11110111011101100101011100001001;
		correct = 32'b00111101100000100100000101010001;
		#400 //-1.2729475e-35 * -4.9963684e+33 = 0.06360114
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100101110110100010010011000;
		b = 32'b01011111000110010110001001101011;
		correct = 32'b01100100011000000110011111111011;
		#400 //1498.1436 * 1.1052514e+19 = 1.6558253e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011110100011001100010001101101;
		b = 32'b01000101110011011001011000101100;
		correct = 32'b11100100111000100001011110111101;
		#400 //-5.071676e+18 * 6578.7715 = -3.3365397e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011101010011101010101111001111;
		b = 32'b00001000000011110100100011101100;
		correct = 32'b00100101111001110101100110101111;
		#400 //9.30764e+17 * 4.3118216e-34 = 4.0132884e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101101111000010011010001110101;
		b = 32'b11001110111101110101101000010111;
		correct = 32'b10111101010110011001100011011110;
		#400 //2.5602834e-11 * -2074938200.0 = -0.0531243
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001010011011001000001000000111;
		b = 32'b11101001100111100110011101011111;
		correct = 32'b10110100100100100101011111000000;
		#400 //1.1387442e-32 * -2.3937304e+25 = -2.7258466e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000111000010111111110100100111;
		b = 32'b01001100011110001110011100101111;
		correct = 32'b11010100000010000001101110101001;
		#400 //-35837.152 * 65248444.0 = -2338318500000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011101101000101011101101111010;
		b = 32'b00101111100101111100110111011001;
		correct = 32'b10001101110000001111111011011110;
		#400 //-4.307489e-21 * 2.7613004e-10 = -1.1894271e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110000011000101000001010110;
		b = 32'b11111011000000100000110110001111;
		correct = 32'b01110001100011101001000001110100;
		#400 //-2.0908387e-06 * -6.752736e+35 = 1.4118881e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010000100110010111111001101010;
		b = 32'b10110010100111011001111101101111;
		correct = 32'b00000011101111010000010000111110;
		#400 //-6.054263e-29 * -1.8349708e-08 = 1.1109396e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101011101111000110000000010101;
		b = 32'b01010110001101011100011111000110;
		correct = 32'b11000010100001011100001011101111;
		#400 //-1.3384872e-12 * 49967406000000.0 = -66.88073
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101000001110001001101111111011;
		b = 32'b10011001010100100010110010010110;
		correct = 32'b11000010000101111001000000011011;
		#400 //3.487171e+24 * -1.08657496e-23 = -37.890728
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010101101011100011100110001011;
		b = 32'b00100011110110000101101011110111;
		correct = 32'b10111010000100110011111001110110;
		#400 //-23945271000000.0 * 2.3457292e-17 = -0.00056169124
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101100111111101110001101101110;
		b = 32'b00011000000110010001100010100101;
		correct = 32'b00000101100110000110111001110110;
		#400 //7.244364e-12 * 1.9787229e-24 = 1.4334588e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010010000001100111111101011;
		b = 32'b10101001101101111100011101001000;
		correct = 32'b00100100100010100110101010111001;
		#400 //-0.0007355201 * -8.161402e-14 = 6.0028755e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111011100000000100101001111;
		b = 32'b01111000111001100011100000001001;
		correct = 32'b11110000110101111101110011100111;
		#400 //-1.4307282e-05 * 3.735515e+34 = -5.3445065e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101100101110100010010110100011;
		b = 32'b10000111101000010000100000011000;
		correct = 32'b00110100111010100010111100011100;
		#400 //-1.8003035e+27 * -2.4229345e-34 = 4.3620173e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010111000000101110101001011010;
		b = 32'b00110001001100011100111010000110;
		correct = 32'b01001000101101011101101101001011;
		#400 //143943040000000.0 * 2.5874285e-09 = 372442.34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110101011000111000100100010101;
		b = 32'b00001011000001011110000110101010;
		correct = 32'b10000000111011011111110110010101;
		#400 //-8.476357e-07 * 2.578464e-32 = -2.185598e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001111010100101011111100101110;
		b = 32'b10100101101110111110101011110110;
		correct = 32'b10110101100110101011001100010100;
		#400 //3535744500.0 * -3.2598545e-16 = -1.1526013e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000011011101010111001000101110;
		b = 32'b00001111001101111110001010100111;
		correct = 32'b10010011001100000100110111101110;
		#400 //-245.44601 * 9.066248e-30 = -2.2252745e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100000000101000000011101011011;
		b = 32'b10000011010100110110111010000111;
		correct = 32'b10100011111101001000001111110010;
		#400 //4.2666377e+19 * -6.2134206e-37 = -2.6510414e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110100010101011110010111110100;
		b = 32'b10010110111100000011010101100100;
		correct = 32'b11001011110010001011010000110001;
		#400 //6.7787063e+31 * -3.8807785e-25 = -26306658.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010101011011011010001110111000;
		b = 32'b00111000001100110100000101010011;
		correct = 32'b00001110001001100110011000011101;
		#400 //4.799092e-26 * 4.2737764e-05 = 2.0510245e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110111011001001100111101001110;
		b = 32'b10110101000101010011100101101111;
		correct = 32'b11101101000001010101111111111110;
		#400 //4.6408138e+33 * -5.55904e-07 = -2.579847e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000010111000101111100111010011;
		b = 32'b01100110110000010001001100110100;
		correct = 32'b01101010001010110010111101011111;
		#400 //113.48794 * 4.558855e+23 = 5.1737505e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000101101010111101111000000011;
		b = 32'b11010111111000111000000110010101;
		correct = 32'b10011110000110001011110011011100;
		#400 //1.6162317e-35 * -500291380000000.0 = -8.085868e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000001011011101011011101110;
		b = 32'b10101100010000011000101111110000;
		correct = 32'b00011101000000110110111000010000;
		#400 //-6.3242467e-10 * -2.750463e-12 = 1.7394607e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011110111100110101101001010101;
		b = 32'b01110101111001111111101101110110;
		correct = 32'b11010101010111001000010110001100;
		#400 //-2.5765986e-20 * 5.8814493e+32 = -15154134000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011000101100001101100100110101;
		b = 32'b10001101000111011010111100100110;
		correct = 32'b10100110010110011101110001101000;
		#400 //1555575500000000.0 * -4.8590187e-31 = -7.5585705e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100111110110101001100101101110;
		b = 32'b01011111110110111111100111110100;
		correct = 32'b11001000001110111101011010110001;
		#400 //-6.0673504e-15 * 3.1701937e+19 = -192346.77
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001110001010110010001111101101;
		b = 32'b11101100011111101001011001000100;
		correct = 32'b00111011001010100011001000011010;
		#400 //-2.1094675e-30 * -1.2311071e+27 = 0.0025969804
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101100100000100000111100101000;
		b = 32'b00110101001010100101011100000101;
		correct = 32'b00100010001011010001010010001101;
		#400 //3.696505e-12 * 6.3456565e-07 = 2.3456751e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110101101101000000010111000011;
		b = 32'b10110001100100000100011110101110;
		correct = 32'b01100111110010101110101101001011;
		#400 //-4.5641128e+32 * -4.1991006e-09 = 1.9165168e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000001100011001100111101100101;
		b = 32'b01111000100011011011110100010010;
		correct = 32'b00111010100110111110110001110011;
		#400 //5.1725474e-38 * 2.2998396e+34 = 0.0011896029
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010010101000111001101001100111;
		b = 32'b10110010010001011000110000110110;
		correct = 32'b11000101011111000111111011011000;
		#400 //351335060000.0 * -1.14987895e-08 = -4039.9277
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010000110011000010001011110110;
		b = 32'b10111110100111100011011111110100;
		correct = 32'b01001111111111000101010001100100;
		#400 //-27398746000.0 * -0.30902064 = 8466778000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100111110010101110100110011000;
		b = 32'b01100000110101001111001101101001;
		correct = 32'b01001001001010001100101001100001;
		#400 //5.6319526e-15 * 1.2275779e+20 = 691366.06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100000011100011101011100001011;
		b = 32'b01011000101101111100110110110001;
		correct = 32'b10111001101011011010001100001001;
		#400 //-2.0484646e-19 * 1616752500000000.0 = -0.00033118602
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101101010000001000110010110101;
		b = 32'b10110100000001000001000110100100;
		correct = 32'b10100001110001101010101110100100;
		#400 //1.094518e-11 * -1.2299876e-07 = -1.3462435e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100110111110110101000000111011;
		b = 32'b10110000000001011111011010000011;
		correct = 32'b00010111100000111000001010101110;
		#400 //-1.743837e-15 * -4.873543e-10 = 8.498665e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101110100001100101100100000000;
		b = 32'b01000010000000000110010000010100;
		correct = 32'b00110001000001101100001000001011;
		#400 //6.109424e-11 * 32.097733 = 1.9609867e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010110010101011011111100111000;
		b = 32'b10000110110010011011101001011111;
		correct = 32'b10011101101010000110111010111111;
		#400 //58754314000000.0 * -7.5881644e-35 = -4.458374e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100010100101001100000001101110;
		b = 32'b00011111000010011100011111111111;
		correct = 32'b01000010001000000001111001100001;
		#400 //1.3719921e+21 * 2.917631e-20 = 40.029667
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111100011011001100101000000110;
		b = 32'b10100100110011010001000110111001;
		correct = 32'b01100001101111011010111000101011;
		#400 //-4.9179183e+36 * -8.89346e-17 = 4.373731e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100111011111100110000110011000;
		b = 32'b10100011011101100100001010100001;
		correct = 32'b00001011011101001011001111111101;
		#400 //-3.5302487e-15 * -1.3349796e-17 = 4.71281e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101110100100010001100001001110;
		b = 32'b01000110001110011000100100101010;
		correct = 32'b11110101010100100101000010011100;
		#400 //-2.2452354e+28 * 11874.291 = -2.6660578e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101101111001111100001011110101;
		b = 32'b01010000010000001110110100000000;
		correct = 32'b11111110101011101010100011000111;
		#400 //-8.965841e+27 * 12947030000.0 = -1.1608101e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000010101011111010000011010100;
		b = 32'b01110001111111110110111011111010;
		correct = 32'b10110101001011110011110101010110;
		#400 //-2.580625e-37 * 2.5296909e+30 = -6.5281836e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010011110010000110001101000110;
		b = 32'b11110111010101010000111001010000;
		correct = 32'b11001011101001101100010111001101;
		#400 //5.058499e-27 * -4.3212872e+33 = -21859226.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111111111010000011111111100000;
		b = 32'b00101000111100001101010110100011;
		correct = 32'b10101001010110100111110110110011;
		#400 //-1.8144493 * 2.6738003e-14 = -4.851475e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111111110110011111100111110000;
		b = 32'b00010110110010000101110010100111;
		correct = 32'b11111111110110011111100111110000;
		#400 //nan * 3.2370215e-25 = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110000010010100100000000111;
		b = 32'b10011010010110101111010111111110;
		correct = 32'b10011000111010101101011010000000;
		#400 //0.13406383 * -4.5280054e-23 = -6.070417e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111000101100101011101110100110;
		b = 32'b10111100001010010101000111010010;
		correct = 32'b01110101011011000110111000000001;
		#400 //-2.9001088e+34 * -0.010334449 = 2.9971025e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011011001011000111010001011;
		b = 32'b10001110110000111010010001010111;
		correct = 32'b00011010101011110110111011110001;
		#400 //-15044235.0 * -4.8229465e-30 = 7.255754e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010101100000111011011001100010;
		b = 32'b01011010111100101011010110101010;
		correct = 32'b01110000111110011011111111000000;
		#400 //18102419000000.0 * 3.4158343e+16 = 6.1834863e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000110010001000101100011010101;
		b = 32'b00110011001110011010110111001000;
		correct = 32'b00111010000011100110100101111011;
		#400 //12566.208 * 4.3231722e-08 = 0.0005432588
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101100100011011000010010111000;
		b = 32'b00000110111011000100101101101101;
		correct = 32'b00110100000000101010000000001100;
		#400 //1.3686823e+27 * 8.888416e-35 = 1.2165418e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110100011100011011101000011111;
		b = 32'b01101011000010011000000001110101;
		correct = 32'b01100000000000011101010111100110;
		#400 //2.2512585e-07 * 1.6622946e+26 = 3.7422547e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111000010011001001110010100;
		b = 32'b11000011100100010001000101011100;
		correct = 32'b11001011000110111110101111010110;
		#400 //35219.58 * -290.13562 = -10218454.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100101001110000110000001111100;
		b = 32'b00100001010001110001011000010111;
		correct = 32'b01000111000011110110001011101001;
		#400 //5.4418453e+22 * 6.745306e-19 = 36706.91
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001110001010100001100011111010;
		b = 32'b01011110001110001100011110110000;
		correct = 32'b00101100111101011000110101000100;
		#400 //2.0966144e-30 * 3.328701e+18 = 6.9790024e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000101101111100110001011000101;
		b = 32'b00111101000101101100101111001001;
		correct = 32'b01000011011000000100101011011010;
		#400 //6092.346 * 0.03681544 = 224.29239
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010000011001111010000101010000;
		b = 32'b10010101111000011111001011000100;
		correct = 32'b10100110110011000111000001101111;
		#400 //15544435000.0 * -9.125979e-26 = -1.4185819e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010110101101111001101010101011;
		b = 32'b00100110000100011110010100100010;
		correct = 32'b00111101010100010100010111100001;
		#400 //100937460000000.0 * 5.0617514e-16 = 0.051092032
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111001111100000001101001100110;
		b = 32'b00101101010011000101101101010100;
		correct = 32'b01100111101111111010101010110001;
		#400 //1.5583583e+35 * 1.1616336e-11 = 1.8102414e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001110011100010010001111010001;
		b = 32'b10110110011010010011111100011100;
		correct = 32'b01000101010110111011010100001011;
		#400 //-1011414100.0 * -3.475644e-06 = 3515.3152
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111011011100111100011111011;
		b = 32'b11101001010100011110101001111101;
		correct = 32'b01100001010000111000101100110100;
		#400 //-1.4214073e-05 * -1.5860802e+25 = 2.254466e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101001101101001001111000111111;
		b = 32'b00111101100110011011100010100011;
		correct = 32'b10100111110110001110100110110001;
		#400 //-8.021057e-14 * 0.0750592 = -6.020541e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110111100001011110101000100011;
		b = 32'b00010011100100111011101011110101;
		correct = 32'b01001011100110101000111001111101;
		#400 //5.4322214e+33 * 3.729237e-27 = 20258042.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110011000110101111000101011100;
		b = 32'b11100110010011110011000001110101;
		correct = 32'b01011001111110101100110011111011;
		#400 //-3.6075434e-08 * -2.4460593e+23 = 8824265300000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100110001100010000010000110001;
		b = 32'b00000100011000010000001101000101;
		correct = 32'b00101011000110111001011011110010;
		#400 //2.0898405e+23 * 2.6450124e-36 = 5.527654e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101110110100001101100010101110;
		b = 32'b01010110101111111001100000100111;
		correct = 32'b01000110000111000100110111001010;
		#400 //9.497235e-11 * 105330105000000.0 = 10003.447
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111000000000111111110111010001;
		b = 32'b11011000101010110011100111010100;
		correct = 32'b11010001001100001001000010110111;
		#400 //3.146922e-05 * -1506118900000000.0 = -47396385000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001110000101011011011100101101;
		b = 32'b10011000010110000110110101011000;
		correct = 32'b10100110111111010010010100000001;
		#400 //627952450.0 * -2.797255e-24 = -1.7565432e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101011110001101100100001100101;
		b = 32'b11010010100011000000010001000000;
		correct = 32'b11111110110110010111000111001000;
		#400 //4.806273e+26 * -300683360000.0 = -1.4451663e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100001111110000110000101110;
		b = 32'b00100111100100011010101101000100;
		correct = 32'b00101100010110010110101101101100;
		#400 //764.1903 * 4.043127e-15 = 3.0897186e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011001101110011100111110111100;
		b = 32'b10110111000111011000011100110001;
		correct = 32'b11010001011001001010110100001101;
		#400 //6537659600000000.0 * -9.389406e-06 = -61384740000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000001010111011111100101001000;
		b = 32'b00010111001101110001011100011111;
		correct = 32'b00011001000111101100000100111111;
		#400 //13.87336 * 5.915967e-25 = 8.207434e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100110100001011011111111011011;
		b = 32'b10101110010010001000010000011101;
		correct = 32'b11010101010100011000010111010010;
		#400 //3.1580693e+23 * -4.5592075e-11 = -14398293000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110101011111101111000100001111;
		b = 32'b00111111110110110100101011011010;
		correct = 32'b00110101110110100110001011000011;
		#400 //9.497316e-07 * 1.7132218 = 1.6271009e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101100000101011110001110011011;
		b = 32'b10110101101100111011110101010110;
		correct = 32'b00100010010100100111101000000010;
		#400 //-2.130052e-12 * -1.3391643e-06 = 2.8524897e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110111100111110001010110100001;
		b = 32'b10101101101010111010010001110000;
		correct = 32'b10100101110101010101001101000100;
		#400 //1.8964349e-05 * -1.9513474e-11 = -3.7006033e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011011011001000111000011100001;
		b = 32'b00100110111101000010110001001100;
		correct = 32'b00000010110110011110001100011110;
		#400 //1.8896191e-22 * 1.6942908e-15 = 3.2015643e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101100000010111000001010101110;
		b = 32'b11110111100011010011011000000110;
		correct = 32'b01100100000110011110100011010101;
		#400 //-1.982563e-12 * -5.7282e+33 = 1.1356517e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000100101001000000011010011011;
		b = 32'b01100010001010101001011101110001;
		correct = 32'b11100111010110101001101011010110;
		#400 //-1312.2064 * 7.8671475e+20 = -1.0323321e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001111010010101101001001110010;
		b = 32'b11011010000101111010111111100101;
		correct = 32'b10101001111100000101101011111001;
		#400 //9.999899e-30 * -1.067403e+16 = -1.0673922e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101010000011101100100001000101;
		b = 32'b10110001101110100100010010100110;
		correct = 32'b11011100010011111100011110011000;
		#400 //4.3153303e+25 * -5.421117e-09 = -2.339391e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011001001000111001110101101001;
		b = 32'b10110000110001010110010000010111;
		correct = 32'b01001010011111000101000000110100;
		#400 //-2878343500000000.0 * -1.4362084e-09 = 4133901.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011001110100000100010110011100;
		b = 32'b10001100000000110010001011101001;
		correct = 32'b00100110010101010110000000001011;
		#400 //-7327916400000000.0 * -1.0102378e-31 = 7.402938e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010000111000110100011001101100;
		b = 32'b01001100010100111010110101101011;
		correct = 32'b01011101101110111110110100000001;
		#400 //30504346000.0 * 55489964.0 = 1.6926851e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100110110100110101000101110001;
		b = 32'b00011100001111011000111111000101;
		correct = 32'b01000011100111000111100111001110;
		#400 //4.9896083e+23 * 6.272067e-22 = 312.9516
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100101000001000100101001110110;
		b = 32'b00100011101000011010001101101100;
		correct = 32'b01001001001001110000111010001111;
		#400 //3.904537e+22 * 1.7524867e-17 = 684264.94
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101011100101101010100010001111;
		b = 32'b10001011101000111110010001001101;
		correct = 32'b10110111110000001110011101011101;
		#400 //3.6426974e+26 * -6.3128825e-32 = -2.299592e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001100110000101010101000110111;
		b = 32'b10001100111110011001011011010010;
		correct = 32'b00011010001111011100101000111111;
		#400 //-102060470.0 * -3.8455296e-31 = 3.9247657e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000100101001111000111000001100;
		b = 32'b00100010001010100111101010001010;
		correct = 32'b10100111010111110010100100010000;
		#400 //-1340.439 * 2.3104168e-18 = -3.0969727e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001101001101101000111101110000;
		b = 32'b10001111010011101010010111001001;
		correct = 32'b10011101000100110101110110100110;
		#400 //191428350.0 * -1.0188513e-29 = -1.9503703e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110110010001101110000111101010;
		b = 32'b10111101111011000110110110111101;
		correct = 32'b01110100101101111010110110000101;
		#400 //-1.008454e+33 * -0.115443684 = 1.1641964e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010111010001011100100011111001;
		b = 32'b00100101101000100011111111011011;
		correct = 32'b00111101011110101011010100000110;
		#400 //217466960000000.0 * 2.814579e-16 = 0.061207794
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101001001001010111000000101000;
		b = 32'b10100111110111101100111011110111;
		correct = 32'b10010001100011111111110100000011;
		#400 //3.673464e-14 * -6.184177e-15 = -2.2717352e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110111110010111010001010110;
		b = 32'b10011100100010001000100010101111;
		correct = 32'b10011100000001010000101011111110;
		#400 //0.4872157 * -9.035057e-22 = -4.4020216e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011000100001101010101111100010;
		b = 32'b00101101000110001010000011101000;
		correct = 32'b10000110001000001001010101100111;
		#400 //-3.4811745e-24 * 8.675928e-12 = -3.020242e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010101010000000101110000111110;
		b = 32'b10110111011010111111000111110000;
		correct = 32'b11001101001100010100101001111000;
		#400 //13218901000000.0 * -1.4063422e-05 = -185902980.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100011011100000101101011000010;
		b = 32'b00111011011100010000111111010010;
		correct = 32'b01011111011000100101010001001011;
		#400 //4.4337584e+21 * 0.0036783111 = 1.6308743e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100011011011110111100100010110;
		b = 32'b10110000000100101010101101100000;
		correct = 32'b10010100000010010011001101011110;
		#400 //1.2981857e-17 * -5.335803e-10 = -6.926863e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010101101001010101111011100100;
		b = 32'b11011100111110110010100010000001;
		correct = 32'b10110011001000100011111000110100;
		#400 //6.679268e-26 * -5.6555803e+17 = -3.7775138e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100101001010110101111101100111;
		b = 32'b00111011101100100010111100100101;
		correct = 32'b10100001011011101000111111001010;
		#400 //-1.4864209e-16 * 0.005437749 = -8.082784e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011111000111100010111011110010;
		b = 32'b11000110000101011001110001011011;
		correct = 32'b01100101101110001110001111011111;
		#400 //-1.1398314e+19 * -9575.089 = 1.0913986e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011011010001100101000101000010;
		b = 32'b11100111100011100001110100001111;
		correct = 32'b01000011010111000010111100101011;
		#400 //-1.6404432e-22 * -1.3422242e+24 = 220.18425
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000000001110010010111100101000;
		b = 32'b00111110101010111011000100011011;
		correct = 32'b10111111011110000110010100111010;
		#400 //-2.8935032 * 0.33533558 = -0.9702946
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011001000111101001001111011111;
		b = 32'b00101101111110011101001110010000;
		correct = 32'b00000111100110101100000011100001;
		#400 //8.198271e-24 * 2.8401975e-11 = 2.3284709e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111101100100110000001000110011;
		b = 32'b00001100110100010001010010010111;
		correct = 32'b01001010111100000010000100111101;
		#400 //2.4425992e+37 * 3.221394e-31 = 7868574.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010101111000011100111001110010;
		b = 32'b01111000000000100111110101111011;
		correct = 32'b01001110011001100011001100001000;
		#400 //9.120249e-26 * 1.0586619e+34 = 965526000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101100010010010001010101101100;
		b = 32'b10101010111111101111110010011100;
		correct = 32'b00010111110010000100100110101101;
		#400 //-2.857571e-12 * -4.5294747e-13 = 1.2943295e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000011110100010001101000010110;
		b = 32'b01100010011001110101111110011000;
		correct = 32'b00100110101111001111110010011111;
		#400 //1.2289905e-36 * 1.0670215e+21 = 1.3113594e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100101110011010100101010010110;
		b = 32'b00111011001000011100110011111001;
		correct = 32'b00100001100000011100000001000111;
		#400 //3.5612373e-16 * 0.0024688824 = 8.792275e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000110010101010101100100101110;
		b = 32'b00100101101101000001011110011111;
		correct = 32'b00101100100101100001011001100100;
		#400 //13654.295 * 3.124103e-16 = 4.2657423e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110011011111010010111100111010;
		b = 32'b01100101010111111010110110101001;
		correct = 32'b01011001010111010011011111100100;
		#400 //5.8949105e-08 * 6.60182e+22 = 3891714000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101100110001001101000100111000;
		b = 32'b01111010010001100011001111101100;
		correct = 32'b01100111100110000110000110111100;
		#400 //5.593883e-12 * 2.5728197e+35 = 1.4392052e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011000101000101110010000110001;
		b = 32'b10110110111000011110101110001010;
		correct = 32'b01010000000011111100000001101110;
		#400 //-1432807700000000.0 * -6.732943e-06 = 9647012000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011101001111011000011010101;
		b = 32'b11010011010000011011001110001110;
		correct = 32'b01011111011111011100001111011100;
		#400 //-21979562.0 * -831941100000.0 = 1.8285701e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111010111011100001110100100100;
		b = 32'b11000001011001100000101100111010;
		correct = 32'b11111100110101011111100010100000;
		#400 //6.1817885e+35 * -14.377741 = -8.8880156e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111110010001000010001111101000;
		b = 32'b10010111000111001010010101100101;
		correct = 32'b00010101111100000000100100110100;
		#400 //-0.19154322 * -5.0615076e-25 = 9.694975e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101000101011110111100011001001;
		b = 32'b00110000101110000000011000110100;
		correct = 32'b10011001111111000100011000100010;
		#400 //-1.9481285e-14 * 1.3389525e-09 = -2.6084516e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100111111101110010100101000001;
		b = 32'b00000101000010100011111111011110;
		correct = 32'b00101101100001010111100111100111;
		#400 //2.334371e+24 * 6.5004594e-36 = 1.5174485e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111111111000000111010101011011;
		b = 32'b01000011000111101011000110111100;
		correct = 32'b01111111111000000111010101011011;
		#400 //nan * 158.69427 = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001100101110101110001111111101;
		b = 32'b01000000011101001100110100111100;
		correct = 32'b10001101101100101011011100100010;
		#400 //-2.8795053e-31 * 3.8250265 = -1.1014185e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010101011110010000011010001001;
		b = 32'b00111111010100100111000110001010;
		correct = 32'b11010101010011001011010111001111;
		#400 //-17112904000000.0 * 0.82204497 = -14067577000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100000101100001100110111000100;
		b = 32'b01110011111011110001101111001011;
		correct = 32'b11010101001001010010001101001100;
		#400 //-2.9951724e-19 * 3.7888265e+31 = -11348189000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000000111111100011110111110011;
		b = 32'b00010010011010101101101110100001;
		correct = 32'b00010011111010010011111010111111;
		#400 //7.945062 * 7.4108094e-28 = 5.887934e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010111011111111101110001001011;
		b = 32'b11111100011010011000000110011010;
		correct = 32'b01010100011010010110000100001000;
		#400 //-8.2672993e-25 * -4.8497352e+36 = 4009421200000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000101011110000110110101101110;
		b = 32'b00011111101001100001110011010100;
		correct = 32'b10100101101000010011001011101111;
		#400 //-3974.8394 * 7.0351427e-20 = -2.7963562e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010010011100010111011100111101;
		b = 32'b11011110011100000010010111110010;
		correct = 32'b00110001011000101000001110010100;
		#400 //-7.6193164e-28 * -4.3261258e+18 = 3.2962122e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000110000100100010010001001011;
		b = 32'b01011100101100111001110101100000;
		correct = 32'b00100011010011010001001001101111;
		#400 //2.7486212e-35 * 4.0445645e+17 = 1.1116976e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111011101101111011011101110111;
		b = 32'b11101010011111011001011111001010;
		correct = 32'b11100110101101011111110100111111;
		#400 //0.0056065875 * -7.664376e+25 = -4.2970995e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001110110010111100001001110100;
		b = 32'b10111011001010011110010000010001;
		correct = 32'b01001010100001110011100011100101;
		#400 //-1709259300.0 * -0.0025923292 = 4430962.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100100100100110100001111001001;
		b = 32'b00011110001000001111100111100000;
		correct = 32'b01000011001110010011010000110111;
		#400 //2.1732447e+22 * 8.5220024e-21 = 185.20396
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111100001010001011000000000;
		b = 32'b10111101101011011110110011010111;
		correct = 32'b11000101101101001101010111111100;
		#400 //68140.0 * -0.08492439 = -5786.748
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000000100000101110111110011001;
		b = 32'b01111100111001011000111101101010;
		correct = 32'b10111101111010101101001101011100;
		#400 //-1.2024566e-38 * 9.535558e+36 = -0.11466095
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011110111001001011110010010101;
		b = 32'b10111110111011001001110111101001;
		correct = 32'b11011110010100110110101011110001;
		#400 //8.2411063e+18 * -0.46214226 = -3.8085634e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110010011100001011011010001110;
		b = 32'b00010111101010101110000110111001;
		correct = 32'b11001010101000001010110101111001;
		#400 //-4.7678142e+30 * 1.1042973e-24 = -5265084.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100000011000100100010111110100;
		b = 32'b01110010111110011011100011001001;
		correct = 32'b01010011110111001011100101011110;
		#400 //1.916609e-19 * 9.8925004e+30 = 1896005500000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110001001101011010111110100001;
		b = 32'b10110100010101010001101110100100;
		correct = 32'b10100110000101110011111010111111;
		#400 //2.64388e-09 * -1.9847226e-07 = -5.2473686e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011001110000101011101111010001;
		b = 32'b10000101000111110010111101110010;
		correct = 32'b10011111011100100010110101111100;
		#400 //6851581500000000.0 * -7.4848584e-36 = -5.1283117e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111001000011100001010110001000;
		b = 32'b01100100110110100101011101100110;
		correct = 32'b01011110011100100101110110101111;
		#400 //0.00013550196 * 3.2221503e+22 = 4.3660768e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111101010001010111100010111;
		b = 32'b11010011101111101001101011101100;
		correct = 32'b01001011111110110011000000010000;
		#400 //-2.0108693e-05 * -1637285900000.0 = 32923680.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100101101101011001110110110110;
		b = 32'b11100100110001010010011110100011;
		correct = 32'b01001011000010111101111001111100;
		#400 //-3.1505364e-16 * -2.9094918e+22 = 9166460.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110010111111101100001010001000;
		b = 32'b11001011011000101101011010110000;
		correct = 32'b01111110111000011011110101100010;
		#400 //-1.0092079e+31 * -14866096.0 = 1.5002982e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110110101011111110101101011100;
		b = 32'b10001011010001000000001001010100;
		correct = 32'b01000010100001101011000111001100;
		#400 //-1.7840344e+33 * -3.7749978e-32 = 67.34726
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101010010011100000000111100110;
		b = 32'b11110110001111100100110111110011;
		correct = 32'b11100001000110010010010000100011;
		#400 //1.8297134e-13 * -9.649584e+32 = -1.7655974e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010010011001010010111001101010;
		b = 32'b10110000100001010111110010010000;
		correct = 32'b10000011011011110000000101000001;
		#400 //7.231687e-28 * -9.712426e-10 = -7.0237227e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111100011101001001100111100001;
		b = 32'b00000111101001111101010010110101;
		correct = 32'b01000100101000000101101110011110;
		#400 //5.080166e+36 * 2.5252385e-34 = 1282.863
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100110000010001110011101100011;
		b = 32'b11110100101101000100101000100011;
		correct = 32'b01011011010000001101010010101110;
		#400 //-4.7498066e-16 * -1.1427211e+32 = 5.427704e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100101001000000111001001001011;
		b = 32'b00100101000001001010000101100110;
		correct = 32'b01001010101001100100000000101101;
		#400 //4.7355436e+22 * 1.1503859e-16 = 5447702.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100011101101001000111000101000;
		b = 32'b11001011100101110101010001111110;
		correct = 32'b11101111110101010111011011100010;
		#400 //6.661315e+21 * -19835132.0 = -1.32128055e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100001100010101000110101010110;
		b = 32'b10011101001001001011101111000011;
		correct = 32'b00111111001100100101000001010100;
		#400 //-3.1947938e+20 * -2.180229e-21 = 0.6965382
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101011010100110100111110101010;
		b = 32'b01000100101001110111000110010011;
		correct = 32'b10110000100010100011011010110111;
		#400 //-7.5072815e-13 * 1339.5492 = -1.0056372e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111111110111011110000011011001;
		b = 32'b00101011001001000111101101011101;
		correct = 32'b10101011100011101000111011110111;
		#400 //-1.7334243 * 5.8435705e-13 = -1.0129388e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010100110000111001010010011010;
		b = 32'b01111110011110000111010111011000;
		correct = 32'b11010011101111011101000111111101;
		#400 //-1.9748581e-26 * 8.2565106e+37 = -1630543700000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100011001100010000010100101001;
		b = 32'b10101011110101001011100011010001;
		correct = 32'b11001111100100110001100000010010;
		#400 //3.2654455e+21 * -1.5114803e-12 = -4935656400.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000010110010001011010011001;
		b = 32'b10011111100100110000010010010110;
		correct = 32'b00010000011110010101011110111011;
		#400 //-7.8976253e-10 * -6.226451e-20 = 4.9174176e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001010011000111001011010000100;
		b = 32'b10010011010100101011100111111010;
		correct = 32'b10011110001110110101011011001110;
		#400 //3728801.0 * -2.659742e-27 = -9.917648e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101101110110011111100000001111;
		b = 32'b01110011011001110110100010011000;
		correct = 32'b01100001110001010000011111100100;
		#400 //2.4780204e-11 * 1.8334076e+31 = 4.5432215e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110101101101000100000101011100;
		b = 32'b01110100101111101101111011000010;
		correct = 32'b01101011000001100110010101011100;
		#400 //1.3430067e-06 * 1.2097833e+32 = 1.6247472e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010010111000001000110101100011;
		b = 32'b11100101110010100101110001010000;
		correct = 32'b10111001001100011000000010001001;
		#400 //1.4171242e-27 * -1.1945261e+23 = -0.00016927918
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101110101001111011100101001111;
		b = 32'b00100011010001101101100100110101;
		correct = 32'b11010010100000100100011110100010;
		#400 //-2.595401e+28 * 1.0779597e-17 = -279773770000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101001110100100110101010100001;
		b = 32'b11010011111011110110100011111010;
		correct = 32'b11111110010001001100011111010101;
		#400 //3.1797245e+25 * -2056516800000.0 = -6.539157e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010011110100111001111100101110;
		b = 32'b01110011000000011111000101110111;
		correct = 32'b01000111010101101101010110100011;
		#400 //5.342085e-27 * 1.0295163e+31 = 54997.637
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100110111101010110101000011111;
		b = 32'b10011000000010001001101001001000;
		correct = 32'b10111111100000101111010001000111;
		#400 //5.794687e+23 * -1.765548e-24 = -1.0230798
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011101111100111110100000100001;
		b = 32'b10111111001100100011101101011100;
		correct = 32'b11011101101010011100111111110101;
		#400 //2.1969167e+18 * -0.69621825 = -1.5295335e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011001101011101000111110111110;
		b = 32'b11010001101010011010111111001001;
		correct = 32'b01101011111001110110100110000011;
		#400 //-6141836500000000.0 * -91099830000.0 = 5.5952026e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011001001010010100101110000010;
		b = 32'b00000111101100100001101100110001;
		correct = 32'b10100001011010111001000011111000;
		#400 //-2978268300000000.0 * 2.6798445e-34 = -7.981296e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111111111100100100111110010001;
		b = 32'b11001000101111111010011001011100;
		correct = 32'b11111111111100100100111110010001;
		#400 //nan * -392498.88 = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000010101110000000001101011101;
		b = 32'b11110111010001100011011101001110;
		correct = 32'b11111010100011100111101001011011;
		#400 //92.00657 * -4.0202988e+33 = -3.698939e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001010100100110110001010011100;
		b = 32'b00110110000011111110001101100101;
		correct = 32'b01000001001001011010110111111111;
		#400 //4829518.0 * 2.1441022e-06 = 10.3549795
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111111001101100110000001110010;
		b = 32'b01010101110000011100011101001011;
		correct = 32'b01010101100010100000110010110000;
		#400 //0.71240914 * 26632713000000.0 = 18973387000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110010101011100000101100110110;
		b = 32'b01011001000101110000011100000100;
		correct = 32'b11001100010011010101101011000100;
		#400 //-2.0261364e-08 * 2656902200000000.0 = -53832464.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101010011110110110001010101000;
		b = 32'b00110000011011100111010111011100;
		correct = 32'b01011011011010100010100101110100;
		#400 //7.597657e+25 * 8.6751384e-10 = 6.5910723e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101011011110000101011011101001;
		b = 32'b00110111011100100000001001011000;
		correct = 32'b10100011011010101100010001101110;
		#400 //-8.822791e-13 * 1.442487e-05 = -1.2726761e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001011110011100101011010101011;
		b = 32'b01100100111000100100011010011111;
		correct = 32'b10110001001101100110000101101111;
		#400 //-7.947872e-32 * 3.3392424e+22 = -2.653987e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000101011010000111101110000111;
		b = 32'b00110101101011101011001111011000;
		correct = 32'b10111011100111101010011101001000;
		#400 //-3719.7205 * 1.3016352e-06 = -0.004841719
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011010111110110110110011110101;
		b = 32'b10101101011010001110011100100101;
		correct = 32'b00001000111001001011110111000010;
		#400 //-1.03987196e-22 * -1.3238998e-11 = 1.3766863e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100100001111110110000100111010;
		b = 32'b11100000110101110100001110001011;
		correct = 32'b01000101101000001110110100100110;
		#400 //-4.1498877e-17 * -1.24091155e+20 = 5149.6436
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001111110011000101101100110111;
		b = 32'b01010111110011000100110110110010;
		correct = 32'b00101000001000110001011010110101;
		#400 //2.0151088e-29 * 449268140000000.0 = 9.0532415e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011011111101101100100111011;
		b = 32'b10000011111101011110110011111011;
		correct = 32'b00001111111101001101000111010000;
		#400 //-16701755.0 * -1.4454214e-36 = 2.4141074e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110011111111000110001010101101;
		b = 32'b01000101001100000000101001010000;
		correct = 32'b00111001101011011000111000000010;
		#400 //1.17526135e-07 * 2816.6445 = 0.00033102935
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111011010001001100100111111111;
		b = 32'b10100000010011000010001001101010;
		correct = 32'b11011100000111001110101101101100;
		#400 //1.02178715e+36 * -1.7290859e-19 = -1.7667578e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100000110001000111010010011010;
		b = 32'b11011010011011001000100111110011;
		correct = 32'b01111011101101011000010101011011;
		#400 //-1.1324887e+20 * -1.6644943e+16 = 1.885021e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101010011110001001000111101100;
		b = 32'b00101101000001111011000111101101;
		correct = 32'b01011000000000111100000110110110;
		#400 //7.5125675e+25 * 7.713369e-12 = 579472000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010101001101110001010010100101;
		b = 32'b01111011010001101011000101001110;
		correct = 32'b01010001000011100001100011000101;
		#400 //3.697284e-26 * 1.03167094e+36 = 38143807000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100011010100110010000100100111;
		b = 32'b00111011001110000101010000011111;
		correct = 32'b00011111000110000000010100110100;
		#400 //1.1445353e-17 * 0.0028126312 = 3.2191556e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011010000011011000101000011110;
		b = 32'b00111101101110001010001110110000;
		correct = 32'b11011000010011000010101110001100;
		#400 //-9959958000000000.0 * 0.09015596 = -897949600000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100000111110100100001001101100;
		b = 32'b10001011101101010010101110001110;
		correct = 32'b10101101001100010001101110001010;
		#400 //1.4426476e+20 * -6.97842e-32 = -1.00674e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111011110101000100110001101000;
		b = 32'b11100101001001001011000011001111;
		correct = 32'b11100001100010001001001110010011;
		#400 //0.006478835 * -4.8608103e+22 = -3.1492388e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000000110101011001110010001100;
		b = 32'b00000100011001000101010010000010;
		correct = 32'b10000101101111101000010111110001;
		#400 //-6.6753597 * 2.6840075e-36 = -1.7916716e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010011101101011010101111010001;
		b = 32'b11001011101101100000110100100000;
		correct = 32'b00100000000000010011000101110111;
		#400 //-4.5860248e-27 * -23861824.0 = 1.0943092e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011111001011011111110111010000;
		b = 32'b11000100000010011110110110001110;
		correct = 32'b01100011101110110111110010010010;
		#400 //-1.2537406e+19 * -551.7118 = 6.917035e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011001101000110110100011010011;
		b = 32'b11010001111011110110010100110100;
		correct = 32'b01101100000110001100111101110111;
		#400 //-5749459600000000.0 * -128524390000.0 = 7.389458e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110110110011001000111011100110;
		b = 32'b11011101001101110100001001111000;
		correct = 32'b11010100100100100110111101000011;
		#400 //6.0963093e-06 * -8.2532806e+17 = -5031455000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010110010000111000101111110111;
		b = 32'b11000000111110110000000110011101;
		correct = 32'b01010111101111111011101101110111;
		#400 //-53751480000000.0 * -7.843947 = 421623750000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010101011001110001001100111110;
		b = 32'b01100001110011111101100000000111;
		correct = 32'b01110111101110111001101110001110;
		#400 //15879364000000.0 * 4.792553e+20 = 7.61027e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111000001101001111001000101100;
		b = 32'b11111111111100111100100010000100;
		correct = 32'b11111111111100111100100010000100;
		#400 //1.4680082e+34 * nan = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001011101001010000001010010011;
		b = 32'b01001010110001111010010001110000;
		correct = 32'b10010111000000001010111011111110;
		#400 //-6.355956e-32 * 6541880.0 = -4.15799e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100011111110111010011001101111;
		b = 32'b01001010011010010110010111010100;
		correct = 32'b11101110111001010110111010010100;
		#400 //-9.284251e+21 * 3823989.0 = -3.5502874e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010001101011010000110010010010;
		b = 32'b11100101101101001110010001000101;
		correct = 32'b00110111111101001000111001001001;
		#400 //-2.7302334e-28 * -1.067796e+23 = 2.9153323e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101001000010011011010110001110;
		b = 32'b11010100010010000010111110100000;
		correct = 32'b10111101110101110101111011101011;
		#400 //3.0577584e-14 * -3439170000000.0 = -0.10516151
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111000110101011010101100000010;
		b = 32'b11011110011000001011110000100100;
		correct = 32'b11010111101110111001001010101001;
		#400 //0.00010188484 * -4.0484645e+18 = -412477150000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100110110010001111010100010000;
		b = 32'b01000110101110000001110100011110;
		correct = 32'b11101110000100001000011011111111;
		#400 //-4.7449695e+23 * 23566.559 = -1.118226e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		$display ("Done.");
		$finish;
	end

endmodule