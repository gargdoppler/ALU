`timescale 1 ns/1 ps
    `include "div.v"


    module alu_tb ();
        reg clock;
        reg [31:0] a, b;
        reg [2:0] op;
        reg [31:0] correct;

        wire [31:0] out;
        wire [49:0] pro;

        alu U1 (
                .clk(clock),
                .A(a),
                .B(b),
                .OpCode(op),
                .O(out)
            );
        /* create a 10Mhz clock */
        always
        #100 clock = ~clock; // every 100 nanoseconds invert
        initial begin
            $dumpfile("alu_tb.vcd");
            $dumpvars(0,clock, a, b, op, out);
            clock = 0;

    op = 3'b010;

		/* Display the operation */
		$display ("Opcode: 010, Operation: DIV");
		/* Test Cases!*/
		a = 32'b11101111100001110100101010111000;
		b = 32'b01011100011010110010000000110110;
		correct = 32'b11010010100100110100110110001100;
		#400 //-8.374161e+28 * 2.6472814e+17 = -316330600000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011001011111001110000111110011;
		b = 32'b11110101001010110010001000010011;
		correct = 32'b00100011101111010010010100100000;
		#400 //-4448758000000000.0 * -2.1693698e+32 = 2.0507144e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111000001001100111010010001101;
		b = 32'b11111011010011100110100100110110;
		correct = 32'b00111100010011100111000111110111;
		#400 //-1.3504456e+34 * -1.0717471e+36 = 0.0126004135
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001000100110110001110001101011;
		b = 32'b00010010011000100110010010010010;
		correct = 32'b11110101101011110110010101100101;
		#400 //-317667.34 * 7.143699e-28 = -4.4468187e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010000100011100111100000000010;
		b = 32'b01101001101010001110111011111111;
		correct = 32'b10100110010101111110010101000011;
		#400 //-19121836000.0 * 2.552852e+25 = -7.4903817e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001100000010001001111111100111;
		b = 32'b11000001010100010001010110011010;
		correct = 32'b00001010001001110100100000000010;
		#400 //-1.0525178e-31 * -13.067774 = 8.054301e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100100000010101010011000110110;
		b = 32'b10011101110000101110001101000100;
		correct = 32'b11000101101101100010000001011110;
		#400 //3.0064766e-17 * -5.158636e-21 = -5828.046
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111100111111010001110000011;
		b = 32'b01111000010100000010001001011000;
		correct = 32'b00001110110001000101101000001110;
		#400 //81735.02 * 1.6885849e+34 = 4.840445e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111011100011111101001101111;
		b = 32'b01110011010100100001110111000101;
		correct = 32'b10000011100100110110100011101110;
		#400 //-1.4423028e-05 * 1.6647127e+31 = -8.663974e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101010001011011001111110100001;
		b = 32'b11110000000110010101101111100110;
		correct = 32'b10111001100100001110100111100111;
		#400 //5.24745e+25 * -1.8984922e+29 = -0.0002764009
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111100100000000110100000001110;
		b = 32'b11001010101011010010010100000100;
		correct = 32'b11110001001111011101101001101011;
		#400 //5.333796e+36 * -5673602.0 = -9.401075e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100011001111000000100000101;
		b = 32'b11010010001101011001000111111110;
		correct = 32'b10110001101000110011001110001010;
		#400 //926.0159 * -194959600000.0 = -4.7497837e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111011100000010001001111001010;
		b = 32'b11111111111101111100111000111011;
		correct = 32'b11111111111101111100111000111011;
		#400 //-0.0039391266 * nan = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110110010000011110111011001101;
		b = 32'b11110011000100101110100101110110;
		correct = 32'b10000010101010001111011111000110;
		#400 //2.8898241e-06 * -1.1639564e+31 = -2.4827596e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101011101110111100101011001111;
		b = 32'b00111011101100001011001111110100;
		correct = 32'b11101111100010000000100001101001;
		#400 //-4.5405373e+26 * 0.005392546 = -8.420026e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000001010010111101011110011001;
		b = 32'b10000110111000111010111100011101;
		correct = 32'b01111001111001010011000101101011;
		#400 //-12.740136 * -8.5645215e-35 = 1.4875479e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000010011000000101010011001110;
		b = 32'b01110100001100100110010000010010;
		correct = 32'b00001101101000001111011010100000;
		#400 //56.082817 * 5.6534333e+31 = 9.920134e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100011000001101000110000111001;
		b = 32'b00101101011110001100011001100010;
		correct = 32'b11110101000010100111010010010010;
		#400 //-2.4819678e+21 * 1.4141218e-11 = -1.7551301e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100100010010100011001111001000;
		b = 32'b10010010000110000101010100001101;
		correct = 32'b11010001101010011110011101111100;
		#400 //4.3845628e-17 * -4.8067576e-28 = -91216640000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011000101111101101110110100011;
		b = 32'b00101010100110101101110000001001;
		correct = 32'b00101101100111011100001011011100;
		#400 //4.9337645e-24 * 2.7508575e-13 = 1.7935368e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100101010010101011101100111;
		b = 32'b00100111011010001010111111010100;
		correct = 32'b01011100101110100100111011010101;
		#400 //1354.7313 * 3.2291784e-15 = 4.1952818e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001000101000001011110111010100;
		b = 32'b01011001101110011010110000010000;
		correct = 32'b10101110010111011010000001010110;
		#400 //-329198.62 * 6532757000000000.0 = -5.039199e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011001011011100100111001101;
		b = 32'b10010110100101111000000011100100;
		correct = 32'b01110100000100101101001111100001;
		#400 //-11389389.0 * -2.4476707e-25 = 4.653154e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010100101010110011101110111111;
		b = 32'b11110101011010001110110000110111;
		correct = 32'b10011110101111000011001011011100;
		#400 //5883534000000.0 * -2.9526462e+32 = -1.992631e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001000110111100001100010001001;
		b = 32'b00011111111110101101001111010111;
		correct = 32'b11101000011000101010110100000100;
		#400 //-454852.28 * 1.0622958e-19 = -4.2817856e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010001010100010100011001001111;
		b = 32'b00010010010011110100010010101000;
		correct = 32'b11111110100000010011110100110110;
		#400 //-56176734000.0 * 6.540231e-28 = -8.589412e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001011000011101001000001000101;
		b = 32'b11001001010001100011100100001011;
		correct = 32'b10000001001110000001111000001101;
		#400 //2.7456742e-32 * -811920.7 = -3.3817023e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100011111010000111100110010011;
		b = 32'b00110101101011010010001010011001;
		correct = 32'b10101101101010111101111011001011;
		#400 //-2.5204979e-17 * 1.2899574e-06 = -1.953939e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010000000100110010010001001110;
		b = 32'b00100011110011001111101111011001;
		correct = 32'b11101011101101111100001100101011;
		#400 //-9874520000.0 * 2.2224386e-17 = -4.4431016e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100010110001100010100101001110;
		b = 32'b10111000011101000010110011111101;
		correct = 32'b01101001110011111100000111100010;
		#400 //-1.8277158e+21 * -5.8216032e-05 = 3.1395404e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000000110001011000111010111100;
		b = 32'b11001010001010011110010000000011;
		correct = 32'b00110110000101001101100001001110;
		#400 //-6.1736736 * -2783488.8 = 2.2179624e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010111111100110000000110001111;
		b = 32'b01100111010001100110000000000110;
		correct = 32'b00110000000111001100110000111101;
		#400 //534376040000000.0 * 9.367999e+23 = 5.704271e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100010001100001100000000111100;
		b = 32'b00001001011101010111111011011001;
		correct = 32'b11011000001110000101000001011100;
		#400 //-2.3954216e-18 * 2.9550446e-33 = -810621100000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001010101011101101111100010110;
		b = 32'b00101010110000001011110101100110;
		correct = 32'b00011111011010000100010001010100;
		#400 //1.6839506e-32 * 3.4237473e-13 = 4.918443e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100101111111100100011010010100;
		b = 32'b01110001101111111001010011010101;
		correct = 32'b10110011101010011110001100110110;
		#400 //-1.5009788e+23 * 1.89733e+30 = -7.911005e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111101101101010010001111111100;
		b = 32'b01101101010110101011101101100100;
		correct = 32'b01001111110101000000000011110000;
		#400 //3.0097139e+37 * 4.230892e+27 = 7113662500.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000011100010000110111000000010;
		b = 32'b00100110010111101111011011100110;
		correct = 32'b00011100100111001010010011010011;
		#400 //8.018618e-37 * 7.735633e-16 = 1.036582e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010011010111000101101110111011;
		b = 32'b01001000110001101011010110001101;
		correct = 32'b00001010000011011111001000001001;
		#400 //2.781313e-27 * 406956.4 = 6.834425e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101011011000111110000010110110;
		b = 32'b00011101110011101100000011101010;
		correct = 32'b11001101000011010001001111110000;
		#400 //-8.095845e-13 * 5.4727214e-21 = -147930880.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100001101111101000100110111101;
		b = 32'b00101011101110000100111111111011;
		correct = 32'b11110101100001000101001011010010;
		#400 //-4.393508e+20 * 1.3096185e-12 = -3.3547997e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111001010001001110001110000100;
		b = 32'b00101001111000111100010100000000;
		correct = 32'b11001110110111010100101010101111;
		#400 //-0.00018776773 * 1.0114999e-13 = -1856329600.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011110101000000110010101010010;
		b = 32'b00111101000111110110000101101100;
		correct = 32'b01100001000000001101000010111010;
		#400 //5.778867e+18 * 0.038911268 = 1.4851397e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001001100111000001100100010110;
		b = 32'b00101011010000010001000001100000;
		correct = 32'b00011101110011101111101111010001;
		#400 //3.7579225e-33 * 6.85901e-13 = 5.478812e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111000001100000000011001001110;
		b = 32'b11011110011101011110011000010111;
		correct = 32'b10011001001101110100000101101000;
		#400 //4.196754e-05 * -4.4297188e+18 = -9.474087e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001011110001101101110001011000;
		b = 32'b00001101000100001111010011110010;
		correct = 32'b10111110001011111001100100101011;
		#400 //-7.659836e-32 * 4.466827e-31 = -0.17148273
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000111110000110010001110000101;
		b = 32'b00111010010000011011100010001110;
		correct = 32'b10001101000000001110111111010100;
		#400 //-2.9361216e-34 * 0.00073898665 = -3.973173e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110101000110011111101100100110;
		b = 32'b11110101100011110000000001100000;
		correct = 32'b10111111000010011101001111101001;
		#400 //1.9519417e+32 * -3.625518e+32 = -0.53838974
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110110110000111110010101010010;
		b = 32'b10111010110110111001011111001110;
		correct = 32'b01111011011001000101111110111100;
		#400 //-1.9866192e+33 * -0.0016753615 = 1.1857854e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111100000111101101000001001101;
		b = 32'b01110011100110100000111001011001;
		correct = 32'b10001000000000111111001111110101;
		#400 //-0.009693217 * 2.4411155e+31 = -3.970815e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010110001110001000100000111;
		b = 32'b01011000011000101110111110110010;
		correct = 32'b10100001111000001000111110011001;
		#400 //-0.001518757 * 998076450000000.0 = -1.521684e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110101001000110110110011000;
		b = 32'b11011110000101001100110111001001;
		correct = 32'b00011000000011010111000010011011;
		#400 //-4.9003393e-06 * -2.6806118e+18 = 1.8280674e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010010101101110110011001011110;
		b = 32'b00101011110001010011010100010110;
		correct = 32'b10100110011011100001001101111101;
		#400 //-1.1574159e-27 * 1.4012426e-12 = -8.259925e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010101001000011010100000011011;
		b = 32'b11001000111011101010100111011001;
		correct = 32'b01001011101011010110011001000000;
		#400 //-11108961000000.0 * -488782.78 = 22727808.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110101011000101010001110110111;
		b = 32'b01000101010000010000100011000010;
		correct = 32'b01101111100101100100100010010100;
		#400 //2.8729971e+32 * 3088.5474 = 9.302099e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000000000100011111000010010110;
		b = 32'b01010110110001101010101110011011;
		correct = 32'b10101000101111000000110110011101;
		#400 //-2.2803092 * 109220170000000.0 = -2.0878097e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010100110110110001101001011100;
		b = 32'b10111011010110001111011110111110;
		correct = 32'b00011001000000010100001001111010;
		#400 //-2.2123746e-26 * -0.003310665 = 6.6825685e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110001001011000001011110010111;
		b = 32'b11010001101000010111001011101100;
		correct = 32'b01011111000010000111000000101100;
		#400 //-8.5215904e+29 * -86677225000.0 = 9.831406e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010111100011010111010101100011;
		b = 32'b01100100001110000111011110111011;
		correct = 32'b00110010110001000101000000011010;
		#400 //311070620000000.0 * 1.3611314e+22 = 2.2853829e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100000011000010010111111111001;
		b = 32'b01010111110000001101110100101101;
		correct = 32'b01001000000101010111001111010010;
		#400 //6.4905847e+19 * 424112350000000.0 = 153039.28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001110110010110000111111010100;
		b = 32'b11110101001011101011000000100011;
		correct = 32'b00011001000101001100101001011100;
		#400 //-1703406100.0 * -2.214434e+32 = 7.692287e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100011010001110101101001101011;
		b = 32'b11010101111101110100110111010101;
		correct = 32'b00001100110011100101110011110010;
		#400 //-1.0806958e-17 * -33989207000000.0 = 3.1795265e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101111001100000010001110101101;
		b = 32'b10100101011110110110010010110001;
		correct = 32'b01001001001100110101110111110110;
		#400 //-1.6019781e-10 * -2.1804895e-16 = 734687.4
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101110101000000101110010111100;
		b = 32'b11100101010100110101110000110011;
		correct = 32'b10001000110000100011101100101111;
		#400 //7.2924305e-11 * -6.2382506e+22 = -1.1689864e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000111111000010111101000011000;
		b = 32'b10000110000111011111011011111101;
		correct = 32'b11000001001101101011010010100000;
		#400 //3.3925998e-34 * -2.9709876e-35 = -11.419098
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111001100111000101101001011111;
		b = 32'b01110101110101101000111011111011;
		correct = 32'b11000011001110101000110101011111;
		#400 //-1.0147891e+35 * 5.4397047e+32 = -186.55223
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000110100011010110010111001111;
		b = 32'b10000010110110101000100001000110;
		correct = 32'b11000011001001011010001111111010;
		#400 //5.31879e-35 * -3.2110438e-37 = -165.64053
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011010110100001101010101101101;
		b = 32'b00110010011100100000101010001001;
		correct = 32'b11100111110111001110000010011111;
		#400 //-2.939073e+16 * 1.4088649e-08 = -2.0861283e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101110011110000111111001110100;
		b = 32'b01110010100100111010010011001111;
		correct = 32'b10111011010101110110111010100101;
		#400 //-1.9226289e+28 * 5.848773e+30 = -0.0032872346
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111110010110010000000010010;
		b = 32'b11010010001110100010001111010001;
		correct = 32'b00100101000010111010111000011001;
		#400 //-2.421442e-05 * -199866200000.0 = 1.2115315e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110110000100111111000001001001;
		b = 32'b11010101010000001011100011000100;
		correct = 32'b10100000010001001000001101000110;
		#400 //2.2044571e-06 * -13243737000000.0 = -1.664528e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010110101000111011010010110010;
		b = 32'b10011101111110111010001100110110;
		correct = 32'b00111000001001101000101100111100;
		#400 //-2.6448105e-25 * -6.6607903e-21 = 3.9707156e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010101101111111010000011111100;
		b = 32'b00100111111110100001101111000111;
		correct = 32'b01101101010001000010010010001111;
		#400 //26337268000000.0 * 6.9419055e-15 = 3.7939537e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001010100110110011110110010011;
		b = 32'b00101101000000110010001110101101;
		correct = 32'b01011101000101111000011000110010;
		#400 //5086921.5 * 7.4544095e-12 = 6.824043e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100101101000010011010001101001;
		b = 32'b01110000011111010100110110111011;
		correct = 32'b00110100101000101110101110110100;
		#400 //9.5158475e+22 * 3.1357471e+29 = 3.0346348e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110111100111000101010011110100;
		b = 32'b01100011010011110110101110000111;
		correct = 32'b11010011110000001111001001001001;
		#400 //-6.341573e+33 * 3.8262242e+21 = -1657397200000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001000011001000100101101011110;
		b = 32'b00100011110000000111000111001111;
		correct = 32'b00100100000101111101100000111101;
		#400 //6.869985e-34 * 2.0864882e-17 = 3.2926067e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111111000111101110011110000100;
		b = 32'b01110010111011000011000000110110;
		correct = 32'b01001011101011000011101110111111;
		#400 //2.1122012e+38 * 9.3563835e+30 = 22574974.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001100010100100001101100011000;
		b = 32'b01111001011111001010110010101110;
		correct = 32'b00010010010101001101111011111101;
		#400 //55077984.0 * 8.1997573e+34 = 6.717026e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101111100101011100101101110001;
		b = 32'b00010101110100011011110100011010;
		correct = 32'b01011001001101101101010110011010;
		#400 //2.7247496e-10 * 8.471278e-26 = 3216456400000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110001110110010100111100100100;
		b = 32'b00111111000111000001111110010011;
		correct = 32'b11110010001100100010101000000001;
		#400 //-2.1521255e+30 * 0.6098568 = -3.528903e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011110101011101101110101010100;
		b = 32'b10100111011000111000000001100010;
		correct = 32'b00110110110001001100010011110110;
		#400 //-1.8514506e-20 * -3.1572175e-15 = 5.8641845e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100100011100010001000110110110;
		b = 32'b01011011000000000010100011101100;
		correct = 32'b01001000111100001100010010111101;
		#400 //1.7787766e+22 * 3.607379e+16 = 493093.9
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111001011000001000000100110110;
		b = 32'b01101111000110101010111111110110;
		correct = 32'b00001001101110011100010110101101;
		#400 //0.0002141044 * 4.7873415e+28 = 4.4723023e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110100110111001100000100001100;
		b = 32'b11111110100110001010000001001101;
		correct = 32'b00110101101110010010001010110000;
		#400 //-1.3991953e+32 * -1.0143749e+38 = 1.379367e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100010110001000000101101111111;
		b = 32'b10111111111100001110010000100101;
		correct = 32'b01100010010100000101011101001000;
		#400 //-1.8081951e+21 * -1.8819624 = 9.60803e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100010000101111110001000011100;
		b = 32'b11011110111100100001100101011110;
		correct = 32'b01000010101000001001101010100111;
		#400 //-7.004378e+20 * -8.722539e+18 = 80.302055
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100001111100001001001000100;
		b = 32'b00101111100010111110111001100001;
		correct = 32'b01010100001011011101110101110001;
		#400 //760.2854 * 2.545333e-10 = 2986978000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010000000010111001110100001100;
		b = 32'b01011101011111111001011001010000;
		correct = 32'b00110010000010111101011011000111;
		#400 //9369301000.0 * 1.1510622e+18 = 8.1397e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111100001000001010000110111000;
		b = 32'b10010110100001101010101110100001;
		correct = 32'b01100101000110001010110011100110;
		#400 //-0.009804182 * -2.175718e-25 = 4.506182e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101000000110011000111110000110;
		b = 32'b10110011100100001100110011111111;
		correct = 32'b01110100000001111011111001010110;
		#400 //-2.9006784e+24 * -6.742811e-08 = 4.301883e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100001000111010100110111010101;
		b = 32'b11001010100001101100110010100111;
		correct = 32'b00010110000101010101111010010100;
		#400 //-5.329668e-19 * -4417107.5 = 1.2065968e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110010110110100000001110000011;
		b = 32'b00011100010011001101001111100011;
		correct = 32'b11010110000010000011110101111011;
		#400 //-2.5380137e-08 * 6.7771795e-22 = -37449410000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101111100011110000000101001100;
		b = 32'b10010110001001100100111000110111;
		correct = 32'b11011000110111000010000111111101;
		#400 //2.601247e-10 * -1.3434053e-25 = -1936308300000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110000011010110000110001011111;
		b = 32'b01100010111000100000011101101101;
		correct = 32'b00001101000001010001101110001110;
		#400 //8.551008e-10 * 2.0847496e+21 = 4.1016957e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010111011001111000011100101011;
		b = 32'b10010101100100001100100001011111;
		correct = 32'b11000001010011001011000010101010;
		#400 //7.481073e-25 * -5.8477267e-26 = -12.793131
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011011111010111111010110100111;
		b = 32'b00100000111101111011111111110011;
		correct = 32'b10111010011100111101000100110001;
		#400 //-3.9036238e-22 * 4.197045e-19 = -0.00093008863
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000010110010000000010001001010;
		b = 32'b01001100010011011001010101110110;
		correct = 32'b00110101111110010001000101010100;
		#400 //100.00838 * 53892570.0 = 1.8556989e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111101101001000000000101011;
		b = 32'b11110110011100000101110111011100;
		correct = 32'b10010000110000000011110110001000;
		#400 //92416.336 * -1.21880365e+33 = -7.582545e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101001011011001000001011111100;
		b = 32'b01000111011000001011010101101100;
		correct = 32'b01100001100001101011100100101001;
		#400 //1.7870316e+25 * 57525.42 = 3.1065074e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001110000100010001110000100011;
		b = 32'b00001000111010011110100000011011;
		correct = 32'b01000100100111101101000011101010;
		#400 //1.7886177e-30 * 1.4077745e-33 = 1270.5286
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111100110100010001101000111;
		b = 32'b11001110110001101101000111111010;
		correct = 32'b10111000010001100111011110010101;
		#400 //78918.555 * -1667824900.0 = -4.7318248e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110101000100110100001110111010;
		b = 32'b00001010110101001111001000100000;
		correct = 32'b01101001101100010000101000000001;
		#400 //5.486032e-07 * 2.0505935e-32 = 2.675339e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010101100100111011101001101;
		b = 32'b00110000001010101111101010001101;
		correct = 32'b11001010000001011001101011110000;
		#400 //-0.0013615877 * 6.2201694e-10 = -2188988.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000001100101100001111011100101;
		b = 32'b00101001101010000101011010101101;
		correct = 32'b01010111011001000100101110010100;
		#400 //18.765085 * 7.4757346e-14 = 251013260000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110010100001100010010100110100;
		b = 32'b10001010000101111000110100000001;
		correct = 32'b11100111111000101001100101000000;
		#400 //1.5616571e-08 * -7.2969054e-33 = -2.1401636e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011001000001101000111111110101;
		b = 32'b01001100110100010000001111001001;
		correct = 32'b01001011101001001100111110100100;
		#400 //2367245600000000.0 * 109583944.0 = 21602120.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010010000110000011011100101011;
		b = 32'b10011110100100110001101110011010;
		correct = 32'b01110011000001000111000110111010;
		#400 //-163440150000.0 * -1.5575646e-20 = 1.0493314e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101000000011010001100001001001;
		b = 32'b01000100010001110101000000011100;
		correct = 32'b01100011001101010011100101011000;
		#400 //2.6652066e+24 * 797.2517 = 3.3429927e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000111011000101000111111000;
		b = 32'b11010010001000100100010111011001;
		correct = 32'b00011110001110100110100001111110;
		#400 //-1.7194557e-09 * -174239140000.0 = 9.8683665e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010111010110111110101111101100;
		b = 32'b11110011110010101110100111110101;
		correct = 32'b10100011000010101011101010000110;
		#400 //241806320000000.0 * -3.215299e+31 = -7.520493e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101101001010101110101010101100;
		b = 32'b11100011010101111010010111111101;
		correct = 32'b10001001010010101110010111110001;
		#400 //9.715489e-12 * -3.9780107e+21 = -2.4422983e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101001001011001011110101001110;
		b = 32'b01110100000111010001111101011011;
		correct = 32'b00110100100011001011100011101111;
		#400 //1.3051825e+25 * 4.97941e+31 = 2.621159e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010000000111111110001001100110;
		b = 32'b01000101010111110000000010001100;
		correct = 32'b10001010001101111000101011101010;
		#400 //-3.1531632e-29 * 3568.0342 = -8.837256e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011111111001101110110011101100;
		b = 32'b11001000010110011111001110110110;
		correct = 32'b10010111000001111001111010000000;
		#400 //9.7800743e-20 * -223182.84 = -4.382091e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010100000000011110100001100111;
		b = 32'b00100010110000001100110110100000;
		correct = 32'b10110000101011000111110100100100;
		#400 //-6.558669e-27 * 5.225942e-18 = -1.2550214e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100010010001110111011101001011;
		b = 32'b11000000011010111001000100100000;
		correct = 32'b01100001010110001100010010001000;
		#400 //-9.198745e+20 * -3.6807327 = 2.4991614e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100010011100100101001100000001;
		b = 32'b00110111010011010011100111110000;
		correct = 32'b01101010100101110010001101010110;
		#400 //1.1175233e+21 * 1.2232442e-05 = 9.135733e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001000101000010101011100001100;
		b = 32'b11111011111110101000111001111100;
		correct = 32'b10001100001001001101100001011110;
		#400 //330424.38 * -2.6019283e+36 = -1.2699211e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111010100001100110101010010110;
		b = 32'b11101001111101111011110000010101;
		correct = 32'b10010000000010101110011010100101;
		#400 //0.0010255154 * -3.7436609e+25 = -2.7393383e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001110001000010100101111000000;
		b = 32'b00111000000010001110100100111001;
		correct = 32'b00010101100101101100110000111010;
		#400 //1.9881254e-30 * 3.2642132e-05 = 6.090673e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010101001001110001100000101;
		b = 32'b01101010111110110101110111110111;
		correct = 32'b10001111001001111110110100000011;
		#400 //-0.0012579864 * 1.5194206e+26 = -8.2793825e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110001100001011110011111011011;
		b = 32'b00110011111101101110110011010010;
		correct = 32'b10111101000010101101001110110011;
		#400 //-3.8971684e-09 * 1.1498345e-07 = -0.0338933
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000110010001000110011110101000;
		b = 32'b00001100010001001010111001000100;
		correct = 32'b11111001011111111010010000011000;
		#400 //-12569.914 * 1.5151732e-31 = -8.2960245e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000000010110100000101010010110;
		b = 32'b01100110100110100011101010010000;
		correct = 32'b10011001001101001111010111011011;
		#400 //-3.406896 * 3.6416236e+23 = -9.355432e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100000011001100101000100110011;
		b = 32'b10110110011010100101000010001000;
		correct = 32'b01101001011110111010000111110110;
		#400 //-6.638441e+19 * -3.4915593e-06 = 1.9012826e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111111110001100100100100010001;
		b = 32'b11011110011100000110011111000010;
		correct = 32'b10100000110100110010010111011010;
		#400 //1.5491048 * -4.330757e+18 = -3.5769838e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110001011011101001111111010111;
		b = 32'b01000100011001110000101100010001;
		correct = 32'b00101100100001000011001100110101;
		#400 //3.4724417e-09 * 924.1729 = 3.7573508e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000011011110000101111100110010;
		b = 32'b10001000101011111001100000110000;
		correct = 32'b11111010001101010000110100011110;
		#400 //248.37186 * -1.05682085e-33 = -2.3501794e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111010000110100000010101111100;
		b = 32'b11000000011001100111110110100111;
		correct = 32'b01111001001010110001000101000110;
		#400 //-1.9993124e+35 * -3.6014192 = 5.551457e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101011010100110100001101011111;
		b = 32'b10111011000111101100001001110000;
		correct = 32'b10101111101010100101010011000100;
		#400 //7.5055755e-13 * -0.002422478 = -3.098305e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111100110000010011000110110101;
		b = 32'b01001101000011100111101101100001;
		correct = 32'b01101111001011011000111011001100;
		#400 //8.024972e+36 * 149403150.0 = 5.3713538e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000011111000000110111110100111;
		b = 32'b10000111101110001010100100011000;
		correct = 32'b00111011100110111001001000101110;
		#400 //-1.3191171e-36 * -2.7784627e-34 = 0.0047476506
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110101010011111111011011010001;
		b = 32'b11001000010011001111000001000001;
		correct = 32'b00101100100000011110001111000110;
		#400 //-7.7472674e-07 * -209857.02 = 3.6916884e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011101111010001001110111011000;
		b = 32'b10011001001111100000001010111010;
		correct = 32'b11000100000111001011001110001010;
		#400 //6.1573095e-21 * -9.8233204e-24 = -626.8053
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011011000011111111011110010001;
		b = 32'b00001111100010001001101101111001;
		correct = 32'b01001011000001101110010101100010;
		#400 //1.1908676e-22 * 1.3470521e-29 = 8840546.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101010010101010110001001110101;
		b = 32'b01011100010110010110000001011110;
		correct = 32'b11001101011110110100110010000100;
		#400 //-6.4491537e+25 * 2.447441e+17 = -263505980.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101110111010001110000000011010;
		b = 32'b00111000110000010010000011000111;
		correct = 32'b00110101100110100101011111101101;
		#400 //1.0589947e-10 * 9.2090624e-05 = 1.1499484e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111101000111011010101001111111;
		b = 32'b11100101100111110100111011001100;
		correct = 32'b10010110111111010101110010011001;
		#400 //0.038492676 * -9.403873e+22 = -4.0932792e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000010000110001001001111001111;
		b = 32'b01111001000000011101001111100000;
		correct = 32'b00001000100101100110110111110011;
		#400 //38.144344 * 4.2131477e+34 = 9.053646e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001100111101111100101110001011;
		b = 32'b01001100011001000100000111001010;
		correct = 32'b01000000000010101111010011010111;
		#400 //129915990.0 * 59836200.0 = 2.1711938
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010110110100010110101111101100;
		b = 32'b10100001110111101111100101101001;
		correct = 32'b11110100011100000111000010100001;
		#400 //115130726000000.0 * -1.5109323e-18 = -7.6198464e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111010100100000111000000000100;
		b = 32'b10110101101101001011010100001011;
		correct = 32'b11000100010011001001111001001111;
		#400 //0.0011019711 * -1.3463736e-06 = -818.4736
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001111010010010101000000000000;
		b = 32'b01111110000011011001101011100000;
		correct = 32'b00010000101101011111100010010100;
		#400 //3377463300.0 * 4.7056326e+37 = 7.177491e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111011101110101110111001001010;
		b = 32'b11000011100111100001100000100100;
		correct = 32'b11110111100101110101100011101000;
		#400 //1.9412006e+36 * -316.1886 = -6.1393755e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010111011101001011101010100011;
		b = 32'b00101111000011110000011011111001;
		correct = 32'b11100111110110110000010000110110;
		#400 //-269082440000000.0 * 1.3008251e-10 = -2.0685519e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001011011110110010111010110111;
		b = 32'b01110100000110010101100001000110;
		correct = 32'b00010110110100011010101011000101;
		#400 //16461495.0 * 4.8596913e+31 = 3.3873542e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011101111111101100011011110;
		b = 32'b00110010111001000110000010111001;
		correct = 32'b11011000010101110000110100001011;
		#400 //-25145788.0 * 2.6586678e-08 = -945804100000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111111000000101010000110111101;
		b = 32'b10101000110111100011010001110101;
		correct = 32'b01010101100101100111111111100010;
		#400 //-0.51028043 * -2.46697e-14 = 20684500000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001000110001110011110011110101;
		b = 32'b11001001010001000010010001100000;
		correct = 32'b10111111000000100000010100111011;
		#400 //408039.66 * -803398.0 = -0.5078923
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100011101111001111001011010101;
		b = 32'b00110000111110001001000010011100;
		correct = 32'b00110010010000101001100110110110;
		#400 //2.0485844e-17 * 1.8085475e-09 = 1.1327236e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101100100010011111000100000110;
		b = 32'b11000011100111101100110001001000;
		correct = 32'b00101000010111100110000010000110;
		#400 //-3.920533e-12 * -317.59595 = 1.2344406e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101101010010010000000001100010;
		b = 32'b11001111000110011111101100111111;
		correct = 32'b00011101101001110001011000011001;
		#400 //-1.1425612e-11 * -2583379700.0 = 4.422738e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111110101110010011000001000011;
		b = 32'b11101000001111110011100000101011;
		correct = 32'b11010101111101111110110100001110;
		#400 //1.2307888e+38 * -3.6120325e+24 = -34074690000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000001111011101111011100110110;
		b = 32'b00110110101011111010001011111000;
		correct = 32'b10001010101011100010011100011110;
		#400 //-8.778212e-38 * 5.2343785e-06 = -1.6770305e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011110010000010111001011100000;
		b = 32'b01011001111010111110101111110100;
		correct = 32'b11000011110100011110100110001111;
		#400 //-3.4848625e+18 * 8300756600000000.0 = -419.82468
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001000101110000000000011001010;
		b = 32'b00111001010010011010100001010001;
		correct = 32'b11001110111010011001011010001110;
		#400 //-376838.3 * 0.00019231557 = -1959479000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101101101010110000101111101011;
		b = 32'b01011001001111100111011010111000;
		correct = 32'b00010011111001011110011011001111;
		#400 //1.9445742e-11 * 3350673600000000.0 = 5.8035322e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111001111111110111001110110010;
		b = 32'b11100010101010101101010001010101;
		correct = 32'b11010110101111110110100000001011;
		#400 //1.6579778e+35 * -1.5756233e+21 = -105226790000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111100001001011101011110101010;
		b = 32'b11101001100100000101100100100001;
		correct = 32'b11010010000100110000111101011000;
		#400 //3.4444127e+36 * -2.1813277e+25 = -157904400000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101000010011000001000011101100;
		b = 32'b11011000100011011111001110100101;
		correct = 32'b00001111001110000000001001101011;
		#400 //-1.1327944e-14 * -1248620700000000.0 = 9.072366e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010101111110110110010000100111;
		b = 32'b10000100101010111100111100011000;
		correct = 32'b11010000101110110100101000110100;
		#400 //1.01536105e-25 * -4.0392092e-36 = -25137619000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100100100011101011000011011011;
		b = 32'b11001001010111001111011111011110;
		correct = 32'b10011010101001010101000000001101;
		#400 //6.188229e-17 * -905085.9 = -6.837173e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101101111001100100111110101110;
		b = 32'b01001111001010100011010110111101;
		correct = 32'b11011110001011010011001001101100;
		#400 //-8.909735e+27 * 2855648500.0 = -3.120039e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010001101000001001011110001001;
		b = 32'b00011010001110010101010010011011;
		correct = 32'b01110110110111011101010000000111;
		#400 //86217140000.0 * 3.8325447e-23 = 2.2496055e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111000111111100010100101001001;
		b = 32'b11001110001101000011010101111010;
		correct = 32'b00101010001101001000011100000100;
		#400 //-0.00012119354 * -755850900.0 = 1.6034055e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100100110010011111111101011010;
		b = 32'b10011111101111100010001001000001;
		correct = 32'b11000100100001111111110010011011;
		#400 //8.760244e-17 * -8.05248e-20 = -1087.8939
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101000010011111011100100010010;
		b = 32'b01011010001011000100111011100101;
		correct = 32'b01001101100110100100111011011011;
		#400 //3.9237752e+24 * 1.212511e+16 = 323607400.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111000010100001100100100001100;
		b = 32'b11010011010001001011110011010110;
		correct = 32'b11100100100001111101011010100000;
		#400 //1.6938679e+34 * -844981700000.0 = -2.0046206e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001111101000100011010001101111;
		b = 32'b11000010000000000001001110110011;
		correct = 32'b01001101001000100001101101111100;
		#400 //-5442690600.0 * -32.019238 = 169981890.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100010101001101010101001101011;
		b = 32'b11010011000100011101101001100101;
		correct = 32'b00001111000100100100001111011001;
		#400 //-4.5174827e-18 * -626434300000.0 = 7.211423e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010001010000100000001001001001;
		b = 32'b11000101001000110110100110010111;
		correct = 32'b11001011100101111111011101001110;
		#400 //52078875000.0 * -2614.5994 = -19918492.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110011110111011011100011101000;
		b = 32'b01000111011111011111001101111111;
		correct = 32'b11101011110111111000001011011000;
		#400 //-3.51333e+31 * 65011.496 = -5.404167e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111001010111110101110110110001;
		b = 32'b11100100100101011011100001110011;
		correct = 32'b01010100001111101111011000100010;
		#400 //-7.2486405e+34 * -2.2094847e+22 = 3280692800000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011000001001001011111111011101;
		b = 32'b10110111000011111000011011011001;
		correct = 32'b11100000100100101110110101000101;
		#400 //724575800000000.0 * -8.554861e-06 = -8.469755e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110101000000100110111010101111;
		b = 32'b11010001000011100100100010111101;
		correct = 32'b01100011011010101010110100010100;
		#400 //-1.6534266e+32 * -38194106000.0 = 4.3290097e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101001110110000110111010001001;
		b = 32'b11010100011010010001000010110011;
		correct = 32'b11010100111011011011101011010000;
		#400 //3.2706246e+25 * -4004030200000.0 = -8168331500000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001101000011111010000101011001;
		b = 32'b11010110000001011000110100100001;
		correct = 32'b10110110100010011010100011111000;
		#400 //150607250.0 * -36710298000000.0 = -4.1025887e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010111001100111110010110101011;
		b = 32'b00100110011101010100100011001010;
		correct = 32'b10110000001110111100000110011010;
		#400 //-5.81279e-25 * 8.51001e-16 = -6.830533e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111101010101001000010010001;
		b = 32'b10111011111001100111111110010001;
		correct = 32'b11001011001111010110111101111110;
		#400 //87329.13 * -0.00703425 = -12414846.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110010010010010000010001000000;
		b = 32'b01110001011110101010011100101001;
		correct = 32'b01000000010011010100111000000101;
		#400 //3.981544e+30 * 1.2411734e+30 = 3.207887
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101111011001010110110101100010;
		b = 32'b01010011000000011110110010101000;
		correct = 32'b01011011111000100000011101101101;
		#400 //7.1004303e+28 * 558021200000.0 = 1.2724302e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110110100111010010110100110011;
		b = 32'b01110100100011110101101101000011;
		correct = 32'b01000001100011000101011011110011;
		#400 //1.5939597e+33 * 9.086297e+31 = 17.542456
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011100111111000001100010001111;
		b = 32'b00001111001110100100100001001100;
		correct = 32'b11001101001011010011100011101101;
		#400 //-1.6682309e-21 * 9.184432e-30 = -181636820.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001111111001011101100110000010;
		b = 32'b01000000100010111100101100100100;
		correct = 32'b10001110110100100111010101101010;
		#400 //-2.2664924e-29 * 4.3685474 = -5.1882063e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011011110110100011000010110000;
		b = 32'b01111001000000011101000001110011;
		correct = 32'b00100010010101110010010000001100;
		#400 //1.22830155e+17 * 4.2127134e+34 = 2.9157016e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001011010110001011011111000111;
		b = 32'b00010100101010111000001000001000;
		correct = 32'b10110110001000011011110110111011;
		#400 //-4.1738346e-32 * 1.7317876e-26 = -2.4101307e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110110000100100111111001001010;
		b = 32'b11000001111111100001011000001101;
		correct = 32'b11110011100100111001100011000101;
		#400 //7.428094e+32 * -31.760767 = -2.338764e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011100001111011110001001011100;
		b = 32'b01100010110001011001100100011010;
		correct = 32'b10111000111101100000000110011011;
		#400 //-2.1379062e+17 * 1.8225204e+21 = -0.00011730493
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101000101000011011011100101011;
		b = 32'b00001001110111101011111001010010;
		correct = 32'b11011110001110011101110000111110;
		#400 //-1.7954027e-14 * 5.3623532e-33 = -3.348162e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100000001011001011111110111100;
		b = 32'b10100101110001011010011110000010;
		correct = 32'b10111001110111111011111000101001;
		#400 //1.4632406e-19 * -3.428756e-16 = -0.00042675555
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011010110000110110110001101001;
		b = 32'b11101010011111001000111110010001;
		correct = 32'b10101111110001100001010110101001;
		#400 //2.750341e+16 * -7.633182e+25 = -3.603138e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110100010010011010001001000;
		b = 32'b10100110010000110101100001010111;
		correct = 32'b01001111101100111100111001101100;
		#400 //-4.0890045e-06 * -6.777394e-16 = 6033299500.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010001000110001101100111000110;
		b = 32'b00101011100001010011101011110100;
		correct = 32'b11100101000100101101100110100011;
		#400 //-41030540000.0 * 9.466581e-13 = -4.334251e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100110001111001010111000110101;
		b = 32'b10110010100001100101111111110111;
		correct = 32'b01110011001100111011101010110101;
		#400 //-2.2275461e+23 * -1.5643293e-08 = 1.4239624e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000101011111001111010011111111;
		b = 32'b11001110111000101001010010100100;
		correct = 32'b00110110000011101110011010001011;
		#400 //-4047.3123 * -1900696000.0 = 2.1293843e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110010110011000110000101011010;
		b = 32'b01110110000001000111110111110111;
		correct = 32'b10111100010001010111001101101111;
		#400 //-8.096337e+30 * 6.718145e+32 = -0.012051447
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111011110011100101110110011011;
		b = 32'b10110101001000101000010111010010;
		correct = 32'b01000110001000101000011110100111;
		#400 //-0.0062977797 * -6.0544437e-07 = 10401.913
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000101111111011110010111100000;
		b = 32'b10011000010111110110000001011100;
		correct = 32'b01101101000100010111110101010101;
		#400 //-8124.7344 * -2.8870724e-24 = 2.8141777e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011001110000111010000100101000;
		b = 32'b11010111010101110011010101000001;
		correct = 32'b00000001111010001011010111100000;
		#400 //-2.0227618e-23 * -236623720000000.0 = 8.548432e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111110001101010111101001101111;
		b = 32'b11111000000010110101000101001100;
		correct = 32'b01000101101001101011110001011001;
		#400 //-6.0306495e+37 * -1.1302784e+34 = 5335.5435
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100111100010010101010010011000;
		b = 32'b00100110110001111101101101100110;
		correct = 32'b11000000001011111110100010100010;
		#400 //-3.8116855e-15 * 1.3867867e-15 = -2.7485738
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110110100011001110010010000111;
		b = 32'b10100101110101010100000111110011;
		correct = 32'b11010000001010010010000110011010;
		#400 //4.198929e-06 * -3.69943e-16 = -11350206000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100010001101111110011101001011;
		b = 32'b10110011100111000000010111101000;
		correct = 32'b00101110000101101101111101110100;
		#400 //-2.492357e-18 * -7.2653904e-08 = 3.4304518e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001010101100100101101011001000;
		b = 32'b11101110001100100111010001001111;
		correct = 32'b00011011111111111101101101100001;
		#400 //-5844324.0 * -1.3807235e+28 = 4.2327982e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101110000010000000000001100100;
		b = 32'b00110111110111001110011110111001;
		correct = 32'b01110101100111011001101110011101;
		#400 //1.0522608e+28 * 2.6333948e-05 = 3.995834e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001110000010101111100010101000;
		b = 32'b00101001111001010011001101101000;
		correct = 32'b00100011100110110011100001110001;
		#400 //1.7129537e-30 * 1.01785605e-13 = 1.6829038e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011110100001111101010111101011;
		b = 32'b00011111011110000011011000010110;
		correct = 32'b00111110100011000001100100011010;
		#400 //1.4382155e-20 * 5.256078e-20 = 0.273629
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011010100111111011000101110011;
		b = 32'b00111001010111010101010100111001;
		correct = 32'b01100000101110001011010010101001;
		#400 //2.2474814e+16 * 0.0002110795 = 1.0647559e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000011110000111011010000010001;
		b = 32'b00101011010111110010111010001011;
		correct = 32'b11010111111000000111101100100000;
		#400 //-391.40677 * 7.9290106e-13 = -493638840000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110101001001100110000110111000;
		b = 32'b00110010010000101000010100010111;
		correct = 32'b11000010010110101111011111101101;
		#400 //-6.198202e-07 * 1.1322547e-08 = -54.742115
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111110001000000000011010110001;
		b = 32'b10101100110001000011111001111010;
		correct = 32'b01010000110100001100000011111001;
		#400 //-0.15627553 * -5.5775913e-12 = 28018460000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110101111101011100001001010010;
		b = 32'b11001100011000000110001110110011;
		correct = 32'b11101001000011000011000010100101;
		#400 //6.2307325e+32 * -58822348.0 = -1.0592458e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111101000110010100100000101100;
		b = 32'b00000001001000010111101000100110;
		correct = 32'b01111011011100110000000111110010;
		#400 //0.037422344 * 2.9658667e-38 = 1.2617676e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100010110111000101010010011100;
		b = 32'b10101110000000010011001101011111;
		correct = 32'b01110100010110100100100001110000;
		#400 //-2.0321902e+21 * -2.937683e-11 = 6.917663e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100111100001111000010001011111;
		b = 32'b10111000101011010111101111101000;
		correct = 32'b10101110010001111111100101110110;
		#400 //3.7613544e-15 * -8.272362e-05 = -4.5468927e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001001100000100010101011110000;
		b = 32'b00010011110010010000001011101001;
		correct = 32'b10110101001001011100011011000001;
		#400 //-3.133674e-33 * 5.0742403e-27 = -6.1756515e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100001110011001011110011001111;
		b = 32'b10111010110111110010110100001111;
		correct = 32'b00100110011010101101100110000011;
		#400 //-1.3873555e-18 * -0.0017026978 = 8.147984e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100101001010101110011110110110;
		b = 32'b01011001100010010100101101010000;
		correct = 32'b10001011000111110101010111101100;
		#400 //-1.4823656e-16 * 4830610000000000.0 = -3.0686927e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100111011111100011111100100110;
		b = 32'b10110100101100010111100100100010;
		correct = 32'b11110010001101110101111100101110;
		#400 //1.200646e+24 * -3.3056955e-07 = -3.6320526e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010000000111100111101001011100;
		b = 32'b01110111111000011000011011000011;
		correct = 32'b00010111101100111110010001001111;
		#400 //10635276000.0 * 9.148438e+33 = 1.1625237e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100000100011011101010100100100;
		b = 32'b10000110011010111001111001011011;
		correct = 32'b11011001100110100001100111110010;
		#400 //2.4027374e-19 * -4.431493e-35 = -5421959000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101001101111001010010000111001;
		b = 32'b00111000001001010001001010100000;
		correct = 32'b01110001000100100100011010001100;
		#400 //2.8506697e+25 * 3.935641e-05 = 7.2432156e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111110100001001101011011000011;
		b = 32'b10000100011100101010010000110010;
		correct = 32'b01111001100011000010011100000001;
		#400 //-0.259451 * -2.8522358e-36 = 9.096408e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101111011001101110010000000100;
		b = 32'b00000010011001100111111101011100;
		correct = 32'b11101100100000000011011111100110;
		#400 //-2.0999386e-10 * 1.6934282e-37 = -1.2400518e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110000101000001100010011110010;
		b = 32'b10110001000111010101111000011010;
		correct = 32'b01111111000000101100010001010100;
		#400 //-3.9804555e+29 * -2.2899997e-09 = 1.7381903e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110101000000100100011110111010;
		b = 32'b01011100001111010000100001010111;
		correct = 32'b01011000001100000110111100001010;
		#400 //1.6514975e+32 * 2.1283176e+17 = 775963800000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110000110011011100101000001101;
		b = 32'b01111011010101001100010110000000;
		correct = 32'b10110100111101111001100101100110;
		#400 //-5.0950953e+29 * 1.1047727e+36 = -4.6118947e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011011100011101100010011001000;
		b = 32'b00010000010011100001011100001000;
		correct = 32'b01001010101100010101100000000100;
		#400 //2.3619096e-22 * 4.064408e-29 = 5811202.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110010110011111101101100111011;
		b = 32'b01001011100010101101001001010111;
		correct = 32'b10100110101111111010011100111010;
		#400 //-2.4197666e-08 * 18195630.0 = -1.3298614e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000110000100010011010001110110;
		b = 32'b10011110101000010010111110010001;
		correct = 32'b10100110111001101001111001100011;
		#400 //2.731001e-35 * -1.7066211e-20 = -1.6002387e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001001111000100000010000000110;
		b = 32'b00111000010100101001011010001110;
		correct = 32'b11010001000010010110000010010011;
		#400 //-1851520.8 * 5.0208117e-05 = -36876923000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011110111010101111111100011;
		b = 32'b11111000010011000001010000010110;
		correct = 32'b00010011000010101101100100101001;
		#400 //-29016006.0 * -1.6556812e+34 = 1.7525117e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100011100001001010101001010101;
		b = 32'b11000100101110110001000110101101;
		correct = 32'b00011110001101011000110010111010;
		#400 //-1.4383607e-17 * -1496.5524 = 9.611162e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001100110101011010110100110101;
		b = 32'b10101101010100111010011000010000;
		correct = 32'b00011111000000010011100111110111;
		#400 //-3.2922091e-31 * -1.2030835e-11 = 2.736476e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101011001100111100111111010111;
		b = 32'b10111101000101001100011101101100;
		correct = 32'b00101101100110101011001011011111;
		#400 //-6.388201e-13 * -0.036322996 = 1.7587208e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110110011010010010111111110001;
		b = 32'b11010101111100010001101000001110;
		correct = 32'b11011111111101111001100010110000;
		#400 //1.1823999e+33 * -33136776000000.0 = -3.5682407e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110111100100000110001011100110;
		b = 32'b11011000011011111011111110010000;
		correct = 32'b10011110100110100010110001111100;
		#400 //1.721219e-05 * -1054424130000000.0 = -1.6323783e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010110010000011111001001111000;
		b = 32'b11111001001000111110011101010101;
		correct = 32'b10011100100101110111011001011110;
		#400 //53311785000000.0 * -5.318977e+34 = -1.0022939e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001000011001101101001001000000;
		b = 32'b00111101001101011000100111110110;
		correct = 32'b00001010101000101011111110001000;
		#400 //6.9460255e-34 * 0.044321023 = 1.5672079e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110111010000100010110110110100;
		b = 32'b01100011001010001011100001010101;
		correct = 32'b00010011100100110101000001101101;
		#400 //1.1573942e-05 * 3.1123355e+21 = 3.7187323e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111000100110000101101101000010;
		b = 32'b01101010100111101101010111110101;
		correct = 32'b01001101011101011000111010100001;
		#400 //2.4721252e+34 * 9.601033e+25 = 257485330.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001100100010011100000011111011;
		b = 32'b10101011010101101001000000100110;
		correct = 32'b00100000101001000101101101101111;
		#400 //-2.1224338e-31 * -7.622812e-13 = 2.7843186e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100010101011010011111100100110;
		b = 32'b01111100010111000010100101110001;
		correct = 32'b10100101110010010111001010101010;
		#400 //-1.5979185e+21 * 4.5725834e+36 = -3.494564e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111011110111011101011110001101;
		b = 32'b11111101001100101000111110100110;
		correct = 32'b00111110000111110000011010001000;
		#400 //-2.303739e+36 * -1.4834278e+37 = 0.15529835
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010001111101111010110110000;
		b = 32'b01010010111010100000011111110100;
		correct = 32'b10100110110100001110001010101110;
		#400 //-0.0007284535 * 502577900000.0 = -1.4494341e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010111100111000011100111000010;
		b = 32'b11101111111110010010111101010100;
		correct = 32'b10100111001000000111111110010011;
		#400 //343543760000000.0 * -1.5423797e+29 = -2.2273619e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010101010111111010101010101100;
		b = 32'b10101100100001111000101010011110;
		correct = 32'b01101000010100110011100011010010;
		#400 //-15370258000000.0 * -3.8523204e-12 = 3.98987e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111111101001011011000101010000;
		b = 32'b01100110111100110110111000110111;
		correct = 32'b00011000001011100011111110000101;
		#400 //1.2944736 * 5.7478408e+23 = 2.2521042e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000011000110001001111111010010;
		b = 32'b11001101010000000010000010000111;
		correct = 32'b00110101010010110101110101001111;
		#400 //-152.6243 * -201459820.0 = 7.5759175e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010000110101111101111001011110;
		b = 32'b10011110110010100010001011100010;
		correct = 32'b11110001100010001011001000100010;
		#400 //28973396000.0 * -2.1402009e-20 = -1.35377e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100100010010010011000111000011;
		b = 32'b01111101101111010101111010001100;
		correct = 32'b10100110000001111111111000101110;
		#400 //-1.4845525e+22 * 3.1464376e+37 = -4.718201e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100010011101011100110010110101;
		b = 32'b00100101110100000110110101011001;
		correct = 32'b11111100000101101111001110001010;
		#400 //-1.13355075e+21 * 3.6156345e-16 = -3.1351364e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100111110001111000101001101000;
		b = 32'b10000110111100001110101000000110;
		correct = 32'b01100000010101000000100100100101;
		#400 //-5.5383656e-15 * -9.062183e-35 = 6.1115136e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110111011011011000101101111111;
		b = 32'b01101100111101000001001001011000;
		correct = 32'b01001001111110010010011101111111;
		#400 //4.817983e+33 * 2.3605162e+27 = 2041071.9
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110010000101001000111100011010;
		b = 32'b00001111011010101101101110001100;
		correct = 32'b11100010001000011110111010111111;
		#400 //-8.647271e-09 * 1.1579374e-29 = -7.467823e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001100011101111001101101110100;
		b = 32'b00110110001101100101101101000110;
		correct = 32'b11010101101011011100110100000110;
		#400 //-64908750.0 * 2.7173242e-06 = -23887010000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101101100011011100100101100110;
		b = 32'b01001000100011011110101000101100;
		correct = 32'b01100100011111111100010011100001;
		#400 //5.485108e+27 * 290641.38 = 1.8872425e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100101001000111000011110100100;
		b = 32'b01111101110110101110101101100111;
		correct = 32'b10100110101111110011101001111011;
		#400 //-4.826549e+22 * 3.6374248e+37 = -1.3269139e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011011011001100111000011110011;
		b = 32'b11000000001010001011001011100100;
		correct = 32'b11011010101011101101100011010100;
		#400 //6.4863434e+16 * -2.6359186 = -2.4607525e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000100110100110110000100011110;
		b = 32'b00111111100010110000000101010110;
		correct = 32'b00000100110000101010010011101010;
		#400 //4.969505e-36 * 1.0859783 = 4.576063e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101110001010000010100010001001;
		b = 32'b00100110010011100001010100100101;
		correct = 32'b11000111010100001110001111000101;
		#400 //-3.823478e-11 * 7.1499263e-16 = -53475.77
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101110000111111101000111011101;
		b = 32'b10111111010101101010111100000111;
		correct = 32'b01101110001111101001001111010001;
		#400 //-1.2365456e+28 * -0.8386082 = 1.4745213e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111001011111001000111111001110;
		b = 32'b01111000101101101001001000111001;
		correct = 32'b01000000001100010001000111110100;
		#400 //8.196097e+34 * 2.9623868e+34 = 2.7667208
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101010101001001110011100010000;
		b = 32'b00111111001101011010100011011000;
		correct = 32'b11101010111010000110001010110111;
		#400 //-9.96775e+25 * 0.7096076 = -1.4046848e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010111100010011110011110010100;
		b = 32'b00110000101100111111010001101100;
		correct = 32'b00100110010001000010111000100111;
		#400 //8.911876e-25 * 1.3093433e-09 = 6.806371e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101110101010111000111011001110;
		b = 32'b10101010000001000001000100010111;
		correct = 32'b01000100001001100100011001101000;
		#400 //-7.801547e-11 * -1.1729884e-13 = 665.1001
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100001111110000110010000000111;
		b = 32'b01000110011000100011001000011100;
		correct = 32'b00011011000011001000111101001011;
		#400 //1.6831611e-18 * 14476.527 = 1.1626829e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011111000010000010001000110111;
		b = 32'b11011000101001111000100111110000;
		correct = 32'b11000101110100000000001101000101;
		#400 //9.809463e+18 * -1473687000000000.0 = -6656.4087
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010011011010001101011001001001;
		b = 32'b01001010100000110010100010010111;
		correct = 32'b00001000011000110011101011011001;
		#400 //2.9388168e-27 * 4297803.5 = 6.8379503e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011100100010110000001111101100;
		b = 32'b01110101100110101100101110101110;
		correct = 32'b00100110011001011110011100010011;
		#400 //3.1303467e+17 * 3.9245353e+32 = 7.97635e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111010010111000111010101101001;
		b = 32'b01010101111100100111000101100111;
		correct = 32'b01100011111010001100100101001101;
		#400 //2.8617167e+35 * 33321110000000.0 = 8.5883e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101000001010101001111011101111;
		b = 32'b10001011000111011100001000001101;
		correct = 32'b11011100100010100110111110111110;
		#400 //9.471359e-15 * -3.0383088e-32 = -3.1173127e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111001000001011100110100000101;
		b = 32'b11110011101001011110001011000011;
		correct = 32'b00000100110011100111110001001110;
		#400 //-0.00012760244 * -2.6285652e+31 = 4.8544523e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010111110010101000111001011011;
		b = 32'b10110100100111110110101000101001;
		correct = 32'b10100010101000101010001111001100;
		#400 //1.308988e-24 * -2.96933e-07 = -4.4083615e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110101110010111100000111110001;
		b = 32'b01010110001010000101101000001001;
		correct = 32'b10011111000110101110101101101000;
		#400 //-1.5181123e-06 * 46276163000000.0 = -3.2805492e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110000110001000111011000101110;
		b = 32'b01101010101110010001111011100110;
		correct = 32'b00000101100001111101011101110010;
		#400 //1.4294466e-09 * 1.11898595e+26 = 1.2774481e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100100010111101000101001110011;
		b = 32'b00100000101100101100011100111110;
		correct = 32'b11000011000111110101010100101011;
		#400 //-4.8255848e-17 * 3.028622e-19 = -159.33269
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001011111100001000000110100000;
		b = 32'b10111001101000011010000010110100;
		correct = 32'b00010001101111100111011110100110;
		#400 //-9.2639675e-32 * -0.00030828046 = 3.0050453e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001010110101010001111010100101;
		b = 32'b11001110111000010000011011101101;
		correct = 32'b00111011011100100111010000100110;
		#400 //-6983506.5 * -1887663700.0 = 0.00369955
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011111101001010011100101000001;
		b = 32'b11001011111001010100010001101001;
		correct = 32'b01010011001110000111110100100111;
		#400 //-2.3811237e+19 * -30050514.0 = 792373700000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100101110010000001101001010100;
		b = 32'b00101000100101111101000000111110;
		correct = 32'b11111100101010001011011011111000;
		#400 //-1.1811987e+23 * 1.6854678e-14 = -7.0081354e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000101101100010001000010010011;
		b = 32'b00101011001101001110001000011001;
		correct = 32'b01011001111110101001100010001000;
		#400 //5666.072 * 6.426262e-13 = 8817057000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101100100101001110110110001001;
		b = 32'b01010101000100011110101110001110;
		correct = 32'b01010111000000101010001101101100;
		#400 //1.440342e+27 * 10027555000000.0 = 143638400000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110000111100010100101100111110;
		b = 32'b10100000101111000011011110000001;
		correct = 32'b11001111101001000001100010010010;
		#400 //1.7556443e-09 * -3.1885168e-19 = -5506147300.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111101010000110101011111100101;
		b = 32'b01011010001010000111100101111001;
		correct = 32'b11100010100101000110100111110001;
		#400 //-1.622849e+37 * 1.1855339e+16 = -1.368876e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101110111100011100110001000111;
		b = 32'b01100000000100011011100001110010;
		correct = 32'b11001110010101000110010011010101;
		#400 //-3.7416422e+28 * 4.200107e+19 = -890844500.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010000000111101010010001000101;
		b = 32'b00000100001011010011111110000011;
		correct = 32'b11001011011010100110101010110110;
		#400 //-3.1286554e-29 * 2.0365215e-36 = -15362742.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011111011011011100001110111111;
		b = 32'b01001111010101000001100110010011;
		correct = 32'b00001111100011110111110100000111;
		#400 //5.034862e-20 * 3558445800.0 = 1.4149047e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001111000000111001011101000111;
		b = 32'b00100010111110110011000000000111;
		correct = 32'b10101011100001100001110010101101;
		#400 //-6.4879336e-30 * 6.8084537e-18 = -9.529232e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011010010011010100010001001101;
		b = 32'b10001100011010110010110100110001;
		correct = 32'b11001101010111110111000100100011;
		#400 //4.244818e-23 * -1.8117341e-31 = -234295860.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011110000011100001000000100011;
		b = 32'b01100111011010000001101110111001;
		correct = 32'b00110110000111001010111110100010;
		#400 //2.55918e+18 * 1.0961004e+24 = 2.3348043e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000010100101011010010110011000;
		b = 32'b11001000010100110100100011000110;
		correct = 32'b00111001101101010101000101011010;
		#400 //-74.823425 * -216355.1 = 0.00034583622
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011111111101100100111000001100;
		b = 32'b00011100010001101010100100100101;
		correct = 32'b11000011000111101011001010100100;
		#400 //-1.0431417e-19 * 6.573132e-22 = -158.69781
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111000001000111010111101000101;
		b = 32'b01010111001010010001111111000111;
		correct = 32'b00100000011101111100010000110000;
		#400 //3.902546e-05 * 185953950000000.0 = 2.0986627e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010101000001111000101101111111;
		b = 32'b11010100101011110111011111001001;
		correct = 32'b10111111110001011100000100001100;
		#400 //9314575000000.0 * -6029031500000.0 = -1.5449538
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001001000101111110001101000000;
		b = 32'b11100100011011001100100110111000;
		correct = 32'b00100100001001000011011000010101;
		#400 //-622132.0 * -1.7471868e+22 = 3.560764e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001110111111101110111001110110;
		b = 32'b00111001010001101010011010011101;
		correct = 32'b10010101001001000100001110100110;
		#400 //-6.2845464e-30 * 0.0001894482 = -3.31729e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010000100110011110100010101001;
		b = 32'b11100111101011111001111010100001;
		correct = 32'b10101000011000000101101000101100;
		#400 //20657293000.0 * -1.6586806e+24 = -1.2454051e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011100111010001001110101011100;
		b = 32'b10011110111001000111110100101010;
		correct = 32'b00111101100000100100111110101111;
		#400 //-1.5393149e-21 * -2.4192206e-20 = 0.06362855
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000110110000011100010101010100;
		b = 32'b10101001011011111111010000011110;
		correct = 32'b00011100110011101011101010010110;
		#400 //-7.288848e-35 * -5.32804e-14 = 1.3680168e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001110011011000011010001100101;
		b = 32'b10110110110001000111110111110110;
		correct = 32'b00010111000110011101111010101110;
		#400 //-2.9114473e-30 * -5.855919e-06 = 4.971803e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101111110110111010100010001010;
		b = 32'b11110111110100100100101111000101;
		correct = 32'b10110111100001011011001011010101;
		#400 //1.3596194e+29 * -8.530618e+33 = -1.593811e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111110000011110001110101110011;
		b = 32'b11101101011100100100011101000010;
		correct = 32'b11010000000101110011100001110010;
		#400 //4.755813e+37 * -4.686345e+27 = -10148235000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000001110111000010111111010001;
		b = 32'b00100011111000001110110011011011;
		correct = 32'b11011101011110101001101101011111;
		#400 //-27.523348 * 2.4386441e-17 = -1.1286332e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000001100111101111100000111011;
		b = 32'b10110110010001001111111101001010;
		correct = 32'b10001010110011101001010100110000;
		#400 //5.8396227e-38 * -2.9354874e-06 = -1.9893197e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110101010001101010010000010111;
		b = 32'b11011010000101010100001001010010;
		correct = 32'b00011010101010100101100100110010;
		#400 //-7.399953e-07 * -1.0503173e+16 = 7.0454455e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011110110111110110001010000111;
		b = 32'b00100000000110011100110011110101;
		correct = 32'b01111110001110011110100101000111;
		#400 //8.048288e+18 * 1.3027419e-19 = 6.1779606e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000101111010011011001001010000;
		b = 32'b11000000010001000000010011111010;
		correct = 32'b01000101000110001001101001011111;
		#400 //-7478.289 * -3.0628037 = 2441.6482
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011111010100011110010100011101;
		b = 32'b00110001010011111010101110010010;
		correct = 32'b11101101100000010101111100001011;
		#400 //-1.5124527e+19 * 3.021999e-09 = -5.004808e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100011001011111110000110011101;
		b = 32'b11010001111101110111010011100101;
		correct = 32'b11010000101101011111010000011101;
		#400 //3.2444374e+21 * -132852260000.0 = -24421394000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010110100101111111011010101000;
		b = 32'b01010000111111111010000111100111;
		correct = 32'b10000101000110000010111010011000;
		#400 //-2.4551028e-25 * 34310404000.0 = -7.1555636e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001110000001111010110000011101;
		b = 32'b10111001011111110100011001001101;
		correct = 32'b00010100000010000000111011001111;
		#400 //-1.6722904e-30 * -0.00024344884 = 6.869166e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111111011010011011010110101110;
		b = 32'b00001101110101001001000111000010;
		correct = 32'b01110001000011001011101011010011;
		#400 //0.91292846 * 1.3100599e-30 = 6.968601e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011010001110001111001110111010;
		b = 32'b01110010100001000111101010011001;
		correct = 32'b00100111001100101011001011111010;
		#400 //1.3014844e+16 * 5.24803e+30 = 2.4799486e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101100100000110111111100001000;
		b = 32'b11111000110010100000010111000100;
		correct = 32'b00110011001001101010000101001110;
		#400 //-1.2717534e+27 * -3.2780028e+34 = 3.8796593e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101100101010111110101101111010;
		b = 32'b10100100111110011000011000001010;
		correct = 32'b11000111001100000110000111001101;
		#400 //4.8862555e-12 * -1.0821361e-16 = -45153.8
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011111100101110001001000001100;
		b = 32'b01011110011010010110111101101110;
		correct = 32'b11000000101001011010110001101101;
		#400 //-2.1771553e+19 * 4.205196e+18 = -5.177298
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011010111111000011011101110111;
		b = 32'b11001001111000001100100101010100;
		correct = 32'b10010000100011111001111010011100;
		#400 //1.04314365e-22 * -1841450.5 = -5.664793e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000010001111011010111010111110;
		b = 32'b00111011111101101011101100000010;
		correct = 32'b01000101110001001100111100010000;
		#400 //47.420647 * 0.0075296173 = 6297.883
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111101100000011011011101000111;
		b = 32'b01010110001011110110110101000010;
		correct = 32'b00100110101111010100101101010010;
		#400 //0.063337855 * 48220950000000.0 = 1.3134925e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110010101001100101001101000001;
		b = 32'b11000010011001001101110010000101;
		correct = 32'b01101111101110100000110001010111;
		#400 //-6.5888204e+30 * -57.21535 = 1.1515826e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011010001111010011010000010001;
		b = 32'b10001100111010010011011000010000;
		correct = 32'b01001100110011111011000100011110;
		#400 //-3.9126343e-23 * -3.5931872e-31 = 108890350.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110010110110000111001010100011;
		b = 32'b11100010111100111000100101000000;
		correct = 32'b11001111011000111000011001111011;
		#400 //8.574381e+30 * -2.2462244e+21 = -3817241300.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101000111011110000010110001101;
		b = 32'b11111010000000101011001011010000;
		correct = 32'b00101110011010100001011000110001;
		#400 //-9.029984e+24 * -1.6965633e+35 = 5.322515e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010111011001010000111010101110;
		b = 32'b11100001110100000011110011111001;
		correct = 32'b00110101000011001100110000010010;
		#400 //-251851210000000.0 * -4.8016454e+20 = 5.2451026e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111001011110111010001111110010;
		b = 32'b01111100000100110000011100001111;
		correct = 32'b10111100110110110001001100001010;
		#400 //-8.166198e+34 * 3.0536432e+36 = -0.026742477
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111110011100001101001000000110;
		b = 32'b11000011011001101000000001111101;
		correct = 32'b11111010100001011011101011011111;
		#400 //8.0026306e+37 * -230.5019 = -3.4718284e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111001011110110001111001011;
		b = 32'b11010111001100000101011111001110;
		correct = 32'b00011111011111101001110111000100;
		#400 //-1.0454048e-05 * -193891160000000.0 = 5.3917093e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110010010111111100010100110010;
		b = 32'b00000111011111100010001001000001;
		correct = 32'b11101010011000010110100111011100;
		#400 //-1.3025145e-08 * 1.9118902e-34 = -6.8127054e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101111011011111100111110111101;
		b = 32'b00011100100101001010110100011010;
		correct = 32'b11010010010011100111011000010100;
		#400 //-2.1810727e-10 * 9.838564e-22 = -221686070000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011001111011001101000010010110;
		b = 32'b10110010011010101000101111111001;
		correct = 32'b00100111000000010011110011011100;
		#400 //-2.4486075e-23 * -1.3652419e-08 = 1.7935338e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011010100011101001101010001000;
		b = 32'b01011000001000111100111100111001;
		correct = 32'b01000001110111101101110000010111;
		#400 //2.0069678e+16 * 720441640000000.0 = 27.857466
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101101000010110001011000001011;
		b = 32'b10110010010011001001011100001111;
		correct = 32'b11111010001011100000100100111001;
		#400 //2.6903165e+27 * -1.190871e-08 = -2.2591168e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011111010111011101111001110111;
		b = 32'b01101000000000010100111111010001;
		correct = 32'b10110110110110111001111001001000;
		#400 //-1.5987347e+19 * 2.4426305e+24 = -6.545135e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110001000101000011001011101011;
		b = 32'b11011101000011001011011000100011;
		correct = 32'b00010011100001101100111110100000;
		#400 //-2.1565778e-09 * -6.337081e+17 = 3.403109e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110011011101001100100011110111;
		b = 32'b11101110100010100000101100000000;
		correct = 32'b10000100011000101111100111101111;
		#400 //5.6993454e-08 * -2.1361115e+28 = -2.6680936e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101111110110101001111101111010;
		b = 32'b00101010000101100001100011100010;
		correct = 32'b01000101001110100110111111111100;
		#400 //3.9767284e-10 * 1.3331309e-13 = 2982.999
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010101011011001011101011111100;
		b = 32'b01000111001001010100010000011111;
		correct = 32'b00001101101101110101100110000111;
		#400 //4.7807325e-26 * 42308.12 = 1.1299799e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111110001000111000111111011011;
		b = 32'b10101010001100011100000110000101;
		correct = 32'b01010011011010111000111011100001;
		#400 //-0.15972845 * -1.5787899e-13 = 1011714400000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101011100011110101101101001101;
		b = 32'b01010101000100100010101100110110;
		correct = 32'b11010101111110110001001100100110;
		#400 //-3.466151e+26 * 10044643000000.0 = -34507458000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000000011000100011010110100110;
		b = 32'b00100001000010100111001001010001;
		correct = 32'b10011110101101011001100100100110;
		#400 //-9.019124e-39 * 4.6907515e-19 = -1.9227461e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010111100110001010100100001010;
		b = 32'b10111110010101101010111000110100;
		correct = 32'b01011000101101100000101011110110;
		#400 //-335703570000000.0 * -0.2096489 = 1601265500000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110010001000110000101001001000;
		b = 32'b11101011111000110101010011101011;
		correct = 32'b11000101101101111001100111001101;
		#400 //3.229343e+30 * -5.4965435e+26 = -5875.225
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001101010111110000010010000111;
		b = 32'b00001010100100011011110001110110;
		correct = 32'b01000010010000111110000001010110;
		#400 //6.872263e-31 * 1.4033883e-32 = 48.969078
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010110000100001011000010100101;
		b = 32'b11011111010000111010101110100000;
		correct = 32'b10110110001111010100110100011100;
		#400 //39772090000000.0 * -1.4099539e+19 = -2.8208078e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101111100001011100010010010110;
		b = 32'b11000000010101111110101110000100;
		correct = 32'b00101110100111101001100100110111;
		#400 //-2.4332242e-10 * -3.3737497 = 7.2122246e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111101110011101110001101111111;
		b = 32'b00101101100100011000000110110000;
		correct = 32'b01001111101101011111111100110101;
		#400 //0.10101985 * 1.6542184e-11 = 6106802700.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111111101000000001110111101011;
		b = 32'b01000100101001110100011101111100;
		correct = 32'b10111010011101010000100111110101;
		#400 //-1.250913 * 1338.2339 = -0.0009347492
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100110111101011110000001110011;
		b = 32'b11000011011011010110101111011000;
		correct = 32'b11100011000001001000111011111111;
		#400 //5.8056007e+23 * -237.42126 = -2.4452742e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110000000010011010010111101011;
		b = 32'b00101110000001010110000010101010;
		correct = 32'b01000001100001000001100100101101;
		#400 //5.0076093e-10 * 3.0326554e-11 = 16.512293
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100011101010011000100101111101;
		b = 32'b10010011000100101111110011011111;
		correct = 32'b01010000000100111010001011101010;
		#400 //-1.8381245e-17 * -1.8552466e-27 = 9907710000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110000101101001100010100000110;
		b = 32'b10100010001010110010100011111011;
		correct = 32'b11001110000001110010111110110111;
		#400 //1.3152721e-09 * -2.3196516e-18 = -567012800.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111111010111111100100001011011;
		b = 32'b10111001101010110110001100000111;
		correct = 32'b01000101001001110010000110111001;
		#400 //-0.87415093 * -0.00032689443 = 2674.1077
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110111100001000111101001101100;
		b = 32'b11111010000110010010111011101010;
		correct = 32'b10111100110111010110010111010000;
		#400 //5.3739547e+33 * -1.9884324e+35 = -0.027026087
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110110100010010110010000101111;
		b = 32'b11001000011110001001110100010101;
		correct = 32'b01101101100011010111100100101001;
		#400 //-1.3933137e+33 * -254580.33 = 5.4729825e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110110110010011010111000010000;
		b = 32'b01010111011111011110110101000100;
		correct = 32'b01011110110010110101001110011000;
		#400 //2.0452775e+33 * 279195490000000.0 = 7.3256106e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000001000110010100001110001111;
		b = 32'b10011111010010110000100101010111;
		correct = 32'b11100001010000010011111001101111;
		#400 //9.578994 * -4.2994648e-20 = -2.2279503e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100010101010100011000101010;
		b = 32'b01110000010101010000100000100011;
		correct = 32'b00010011100000000010010101000101;
		#400 //853.0963 * 2.6372058e+29 = 3.2348493e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000001001000101111001110110010;
		b = 32'b01010001011100000110000111101111;
		correct = 32'b10101111001011011000100111101110;
		#400 //-10.184496 * 64527200000.0 = -1.5783261e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011110110110010101111101101000;
		b = 32'b11001001100011001010011010001011;
		correct = 32'b11010100110001011101001001001101;
		#400 //7.831676e+18 * -1152209.4 = -6797094600000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100010110100100100011010101100;
		b = 32'b11001010010001100100011111010111;
		correct = 32'b10011000000001111011111001100000;
		#400 //5.699544e-18 * -3248629.8 = -1.7544456e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110011011001110000101100101011;
		b = 32'b01000010111010100001110000110101;
		correct = 32'b11101111111111001010010110001111;
		#400 //-1.8305162e+31 * 117.05509 = -1.5638074e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101100000111000001010111110010;
		b = 32'b11100001001110011000110011000101;
		correct = 32'b00001010010101110101100101001011;
		#400 //-2.2181115e-12 * -2.1392445e+20 = 1.03686676e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000001111001011101111100011010;
		b = 32'b11000111111101011111101101111010;
		correct = 32'b00111001011011110011101110101001;
		#400 //-28.733936 * -125942.95 = 0.00022815041
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110001100010110011011100010000;
		b = 32'b01101001111010111001100100001010;
		correct = 32'b11000111000101110100010101010001;
		#400 //-1.3787195e+30 * 3.5602534e+25 = -38725.316
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000001101000001010011101010001;
		b = 32'b11110111110010011101111110101111;
		correct = 32'b10001001010010111011101001010111;
		#400 //20.081697 * -8.188973e+33 = -2.4522853e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000110010110011110011010110110;
		b = 32'b10011010001101001100001000000100;
		correct = 32'b11101011100110100100110101100011;
		#400 //13945.678 * -3.7379852e-23 = -3.7308005e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010111111011101000101000010101;
		b = 32'b11001111010101001011110011010010;
		correct = 32'b01001000000011111000011001000001;
		#400 //-524553650000000.0 * -3569144300.0 = 146969.02
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001100101101100100111011101010;
		b = 32'b11100001100110110000100010010101;
		correct = 32'b10101010100101101000010011001111;
		#400 //95582030.0 * -3.5748297e+20 = -2.6737507e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000101000111011001111110100000;
		b = 32'b00001101110110011110110110000000;
		correct = 32'b11110110101110010010100100011100;
		#400 //-2521.9766 * 1.3430834e-30 = -1.8777514e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110010101110010011000111100110;
		b = 32'b01010101100001100000111101011011;
		correct = 32'b10011100101100001101001011001110;
		#400 //-2.1559526e-08 * 18425064000000.0 = -1.1701195e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001010001101001000110011111101;
		b = 32'b11001010101101101011101010100111;
		correct = 32'b10111110111111001111001010111001;
		#400 //2958143.2 * -5987667.5 = -0.49403933
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100100000110100001101101011011;
		b = 32'b01010001110110110000001011011001;
		correct = 32'b11010001101101000010001001010000;
		#400 //-1.1371079e+22 * 117580700000.0 = -96708720000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000011000110100110100011101000;
		b = 32'b00000010001100000011110111110110;
		correct = 32'b01000000011000000100100110100001;
		#400 //4.537696e-37 * 1.294822e-37 = 3.504494
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011000101000110001100100001010;
		b = 32'b11100010001001000110010110110100;
		correct = 32'b00110101111111011111100111111001;
		#400 //-1434623500000000.0 * -7.581486e+20 = 1.892272e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101010011000100010101001100010;
		b = 32'b10110000111100110011011110110100;
		correct = 32'b00111000111011100000110101000010;
		#400 //-2.0087537e-13 * -1.7696409e-09 = 0.00011351194
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011010001101001010101111011110;
		b = 32'b11010101100000000001101111000011;
		correct = 32'b01000100001101001000010010110111;
		#400 //-1.2713616e+16 * -17607090000000.0 = 722.07367
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110101011100011001101100101010;
		b = 32'b01011100000111100110010101100010;
		correct = 32'b00011000110000110011110111111110;
		#400 //9.000529e-07 * 1.7833807e+17 = 5.0468915e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000010001101010100111101100011;
		b = 32'b00001000010100111011110000001110;
		correct = 32'b10111001010110110011011100000111;
		#400 //-1.3320563e-37 * 6.371656e-34 = -0.00020905967
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001110110011111010010001111100;
		b = 32'b01000100000010100010000011110111;
		correct = 32'b11001010010000000110101010011010;
		#400 //-1741831700.0 * 552.5151 = -3152550.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111011110101010010011110000110;
		b = 32'b10010110011010111010000001100101;
		correct = 32'b11100100111001111001010110110101;
		#400 //0.0065049557 * -1.903376e-25 = -3.4175883e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011101111001010010101100100000;
		b = 32'b11010101100000100111110010001001;
		correct = 32'b00000111111000001100110100110100;
		#400 //-6.0660385e-21 * -17933923000000.0 = 3.3824382e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000001011101000111011110110100;
		b = 32'b00000001011011101101010101000001;
		correct = 32'b10111111100000110000010100010001;
		#400 //-4.4901605e-38 * 4.3866698e-38 = -1.0235921
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100010011111011101110011010110;
		b = 32'b10100000000101100111000010101111;
		correct = 32'b01000001110101111111111011100001;
		#400 //-3.4404803e-18 * -1.2742778e-19 = 26.999453
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001100110001010011111111011011;
		b = 32'b00110011101110101001000001010101;
		correct = 32'b11011000100001110101010011010010;
		#400 //-103415510.0 * 8.687554e-08 = -1190387000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110111110010110001001011111100;
		b = 32'b00111100101011010100100010001101;
		correct = 32'b11111010100101100000000101110011;
		#400 //-8.2376665e+33 * 0.021152759 = -3.8943696e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000111101010100101111001111101;
		b = 32'b10111100111101111110010111000111;
		correct = 32'b01001010001011111111000000000011;
		#400 //-87228.98 * -0.030260934 = 2882560.8
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010101111100100100110111001101;
		b = 32'b01100110101010001100111010000101;
		correct = 32'b10101110101101111011101011110010;
		#400 //-33301996000000.0 * 3.985836e+23 = -8.355085e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000010111011110010101100011110;
		b = 32'b10101001001100101111110100110010;
		correct = 32'b00011001001010110000100100110011;
		#400 //-3.5142642e-37 * -3.974355e-14 = 8.8423506e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001101000001101101111000000101;
		b = 32'b11010100000100100111101001011001;
		correct = 32'b00111000011010111011010101000000;
		#400 //-141418580.0 * -2516471500000.0 = 5.619717e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011000001110001010111101011100;
		b = 32'b00000010101101000110010001001001;
		correct = 32'b01010101000000110000101111011110;
		#400 //2.3869976e-24 * 2.6506184e-37 = 9005437000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000010000011011100001101111101;
		b = 32'b11101101101111110011011011000110;
		correct = 32'b00010011101111011100101110010001;
		#400 //-35.440907 * -7.397232e+27 = 4.791104e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011010101111001101010101101011;
		b = 32'b01001000101110110011110000001000;
		correct = 32'b01010001100000010001011111011111;
		#400 //2.6575976e+16 * 383456.25 = 69306410000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001000100110101110011111001010;
		b = 32'b10010000111110110000010010010001;
		correct = 32'b00110111000111011111101011011111;
		#400 //-9.323031e-34 * -9.900908e-29 = 9.41634e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101000110001010000010110100011;
		b = 32'b01100101101110000101110001001011;
		correct = 32'b00000010100010001100101001110000;
		#400 //2.1873838e-14 * 1.0882724e+23 = 2.0099597e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110110111101100100111100010011;
		b = 32'b01010100100111010000101000111110;
		correct = 32'b11100001110010001100001011011101;
		#400 //-2.4978688e+33 * 5395853600000.0 = -4.6292377e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010010011100001000011010110101;
		b = 32'b10101010111011110001011000001011;
		correct = 32'b01100111000000001100010101011111;
		#400 //-258263040000.0 * -4.2470224e-13 = 6.0810376e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010001011100001110100001010111;
		b = 32'b10111110000101101111011101001011;
		correct = 32'b11010010110011000100001001010001;
		#400 //64668135000.0 * -0.14742772 = -438642970000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111111110001100000000010110000;
		b = 32'b00001100100001000010000010010101;
		correct = 32'b11111111110001100000000010110000;
		#400 //nan * 2.035743e-31 = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011011100100010100001100000011;
		b = 32'b11011100110011000011111101101011;
		correct = 32'b10111110001101100001000101110100;
		#400 //8.17751e+16 * -4.59925e+17 = -0.17780095
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111110001100110011010111011100;
		b = 32'b11111011101100000111100100100111;
		correct = 32'b11000010000000011111110000111101;
		#400 //5.9552866e+37 * -1.832603e+36 = -32.496326
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010100010011101111101110010101;
		b = 32'b10010100000100101000001010010111;
		correct = 32'b10111111101101001101010100011111;
		#400 //1.0449958e-26 * -7.3968706e-27 = -1.4127539
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001100111110110011000100101001;
		b = 32'b10011110010101000010001010010010;
		correct = 32'b11101110000101111001000100001011;
		#400 //131696970.0 * -1.12303355e-20 = -1.1726896e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000111011100101000011101010111;
		b = 32'b00000001100110000011111000111010;
		correct = 32'b11000101010010111110100010011001;
		#400 //-1.8245829e-34 * 5.592527e-38 = -3262.5374
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110101101011011000010110000111;
		b = 32'b00011100111000100100011110001001;
		correct = 32'b01011000010001000101000000001101;
		#400 //1.2928366e-06 * 1.4973917e-21 = 863392400000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001010100100100000000010011001;
		b = 32'b00001101000010001010010001110101;
		correct = 32'b10111101000010001100010010010111;
		#400 //-1.4059513e-32 * 4.2106194e-31 = -0.033390608
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000101010001111101111101111001;
		b = 32'b00011110100111111110011100100111;
		correct = 32'b01100110000111111111111011010011;
		#400 //3197.967 * 1.6930382e-20 = 1.8888924e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100100110001110001100010011110;
		b = 32'b00110111111110111101110011110110;
		correct = 32'b00101100010010100101110111001000;
		#400 //8.6344196e-17 * 3.0024425e-05 = 2.8757986e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011001101001111011111001111001;
		b = 32'b10100110101000100010001100001101;
		correct = 32'b11110010100001000110110100110100;
		#400 //5901968500000000.0 * -1.1250509e-15 = -5.245957e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001010100110000011011010110100;
		b = 32'b00010100101101001010111111100100;
		correct = 32'b10110101010101111010100010010011;
		#400 //-1.4657645e-32 * 1.8244732e-26 = -8.033905e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000010000111100110010100101000;
		b = 32'b11000011111100110011101000111101;
		correct = 32'b10111101101001101011011001111111;
		#400 //39.598785 * -486.455 = -0.08140277
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011010001111011110100010111010;
		b = 32'b00110000110011110111110001100111;
		correct = 32'b11101000111010100101000000110111;
		#400 //-1.3363664e+16 * 1.509659e-09 = -8.8521077e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001011000010001100111100100000;
		b = 32'b00101100101010110100010100101000;
		correct = 32'b10011101110011000111110110010101;
		#400 //-2.634847e-32 * 4.86779e-12 = -5.41282e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001110100110101010101111111110;
		b = 32'b00101000000010110100110001101100;
		correct = 32'b00100110000011100010000001011011;
		#400 //3.8129554e-30 * 7.732621e-15 = 4.9309997e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100101100010010000111110110111;
		b = 32'b10101101110111101011011110010100;
		correct = 32'b11110111000111011000101100111011;
		#400 //8.090676e+22 * -2.5320003e-11 = -3.1953693e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111111011111001000000001101;
		b = 32'b00110010101101011010110010010111;
		correct = 32'b11000100101010001100100100101100;
		#400 //-2.8558099e-05 * 2.1149658e-08 = -1350.2866
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110100011010110111000001100000;
		b = 32'b01101101110000110011110101110011;
		correct = 32'b11000110000110100101101011000100;
		#400 //-7.4613586e+31 * 7.552983e+27 = -9878.691
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110100111011111111010000001001;
		b = 32'b00000010111111100001110111001100;
		correct = 32'b11110001011100011011101101011101;
		#400 //-4.4694778e-07 * 3.7339048e-37 = -1.1969983e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111001100000100101100101110110;
		b = 32'b11101110010100101111001011001100;
		correct = 32'b01001010100111100011000000010010;
		#400 //-8.460163e+34 * -1.6321344e+28 = 5183497.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000000011010011111000000111000;
		b = 32'b01110011111011000010001010110100;
		correct = 32'b00001011111111011001111000110011;
		#400 //3.6552868 * 3.7417173e+31 = 9.7690087e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101010100100001101001011100011;
		b = 32'b11011100111111111111110110010001;
		correct = 32'b01001101000100001101010001000011;
		#400 //-8.75406e+25 * -5.7643935e+17 = 151864370.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110110001010010011110010100100;
		b = 32'b11111001110011011110111011110101;
		correct = 32'b10111011110100100110000110111100;
		#400 //8.581329e+32 * -1.33658435e+35 = -0.0064203423
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110111111011011001100000110110;
		b = 32'b00111010111100010001011110111001;
		correct = 32'b11111100011111000100100100011110;
		#400 //-9.637981e+33 * 0.0018393911 = -5.2397672e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010101100011110011011010100010;
		b = 32'b01000110111001100101011111010000;
		correct = 32'b11001110000111110010101001010110;
		#400 //-19683101000000.0 * 29483.906 = -667588000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011111111100011100000100111100;
		b = 32'b11011101100101000110100011011111;
		correct = 32'b00000001110100001000001000010100;
		#400 //-1.0238715e-19 * -1.3367553e+18 = 7.6593786e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101000010111010100001000111110;
		b = 32'b00101000011111110100110111111110;
		correct = 32'b11111111010111011101110010000011;
		#400 //-4.1794598e+24 * 1.41722554e-14 = -2.9490435e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100111000010111000100010001011;
		b = 32'b01011010001001111100010010111000;
		correct = 32'b01001100010101001110101001101111;
		#400 //6.589277e+23 * 1.1805654e+16 = 55814588.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110000001011101110011100010000;
		b = 32'b11100101111001000101111010111100;
		correct = 32'b10001001110001000001000001001010;
		#400 //6.362919e-10 * -1.3480589e+23 = -4.72006e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101001010101010001111100000101;
		b = 32'b01010101010011010111111110100110;
		correct = 32'b01010011100001001011111101110110;
		#400 //1.610298e+25 * 14121758000000.0 = 1140295700000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100011110000011101110011010111;
		b = 32'b01010110010110101000011000101100;
		correct = 32'b00001100111000110001101111110110;
		#400 //2.1018631e-17 * 60067450000000.0 = 3.4991716e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000011010000011000100100000100;
		b = 32'b11010101110001001101111100101001;
		correct = 32'b00101100111110111010100101010011;
		#400 //-193.53522 * -27057843000000.0 = 7.152648e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010000000010011001100000011000;
		b = 32'b11110011110000111001111011001101;
		correct = 32'b00011011101101000001000001000111;
		#400 //-9233785000.0 * -3.0997276e+31 = 2.978902e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101111101001000000010100110111;
		b = 32'b11000111011010110000110011001100;
		correct = 32'b11100111101100101010001110110111;
		#400 //1.0152369e+29 * -60172.797 = -1.6872025e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001100011111100011111000101000;
		b = 32'b00010100110111010100111100101110;
		correct = 32'b01110111000100110000110001000110;
		#400 //66648224.0 * 2.2346528e-26 = 2.9824866e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110000010001011111010110001110;
		b = 32'b10111100111101011000010100100100;
		correct = 32'b01110010110011100110100010110100;
		#400 //-2.4506162e+29 * -0.029970713 = 8.176703e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011101101110001011010001011000;
		b = 32'b11001011011111001111101110100010;
		correct = 32'b11010001101110101110100001000001;
		#400 //1.66367e+18 * -16579490.0 = -100345060000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010111111000001100100101111000;
		b = 32'b10111011000101110011111111010000;
		correct = 32'b11011100001111100011101111011111;
		#400 //494311800000000.0 * -0.0023078807 = -2.141843e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110011011100110011011101010101;
		b = 32'b10010101101000100011000101100010;
		correct = 32'b01011101001111111111000100110101;
		#400 //-5.662817e-08 * -6.550919e-26 = 8.644309e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010100000111100011011101100111;
		b = 32'b01111100011101101100001010000111;
		correct = 32'b10010111001001000010010000010110;
		#400 //-2718137300000.0 * 5.125002e+36 = -5.3036805e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110010100110000000001100101010;
		b = 32'b00100000110010010100100111111001;
		correct = 32'b01010001010000010101010001110001;
		#400 //1.7696568e-08 * 3.4099675e-19 = 51896586000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001100101011110111101110111110;
		b = 32'b01011001000100101000001001101011;
		correct = 32'b00110011000110010101000000111111;
		#400 //92003820.0 * 2577421400000000.0 = 3.5696072e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001010010101101010101111001111;
		b = 32'b01100110011100100111000101101000;
		correct = 32'b00100011011000101010110011011000;
		#400 //3517171.8 * 2.8622617e+23 = 1.2288086e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000001101011000101001001100000;
		b = 32'b00011010001100111011000001110000;
		correct = 32'b01100110111101011000000011110110;
		#400 //21.540222 * 3.7158857e-23 = 5.7967935e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110100100100101010011100101100;
		b = 32'b11000001110011111111101100001101;
		correct = 32'b10110010001101001000001101000111;
		#400 //2.7316253e-07 * -25.997583 = -1.0507228e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111011010011111010110000101101;
		b = 32'b10011100000000000101010111000110;
		correct = 32'b01011110110011110010000101100000;
		#400 //-0.0031688318 * -4.2462507e-22 = 7.462658e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001111110101001010011100110110;
		b = 32'b10100001010100110010110001110101;
		correct = 32'b11101110000000001110010110010100;
		#400 //7135456000.0 * -7.154842e-19 = -9.972906e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111001100010101100111110001000;
		b = 32'b01010000100001001000100100000111;
		correct = 32'b10101000100001100000111110001000;
		#400 //-0.00026476034 * 17788582000.0 = -1.4883724e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100000100000000001000101110101;
		b = 32'b01001111110001111001001100101011;
		correct = 32'b10010000001001000100011011000111;
		#400 //-2.1695596e-19 * 6696621600.0 = -3.2397822e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101111011011101100011000110001;
		b = 32'b00000010011100110001100100100100;
		correct = 32'b01101100011110110111001001001101;
		#400 //2.1716386e-10 * 1.7860035e-37 = 1.2159206e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100101100110010111010101100101;
		b = 32'b01100000000110000000111110111100;
		correct = 32'b01000101000000010010110100010001;
		#400 //9.058595e+22 * 4.3828733e+19 = 2066.8167
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011010010110101011110111010100;
		b = 32'b11111000111011110110011110010000;
		correct = 32'b10100000111010011110011110010101;
		#400 //1.5392566e+16 * -3.8845608e+34 = -3.9624983e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100111001011110111101111001111;
		b = 32'b01010010101011001000111101111101;
		correct = 32'b11010100000000100010101100010101;
		#400 //-8.28698e+23 * 370570850000.0 = -2236274200000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100100000011110100010001111010;
		b = 32'b11011001101110101101101100101001;
		correct = 32'b11001001110001000100100000101101;
		#400 //1.0571275e+22 * -6574414400000000.0 = -1607941.6
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010111110111111110000010000100;
		b = 32'b00111011100100001111101000101001;
		correct = 32'b11011011110001011010100100010100;
		#400 //-492310760000000.0 * 0.0044243527 = -1.1127295e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101101111010110000101111011101;
		b = 32'b01101100101001110100100100011010;
		correct = 32'b00000000101100111101100100000111;
		#400 //2.6721675e-11 * 1.6178866e+27 = 1.6516409e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011110110010011101001111010110;
		b = 32'b00100110000100001010010101011010;
		correct = 32'b01111000001100101001100111100010;
		#400 //7.2716015e+18 * 5.018413e-16 = 1.4489843e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111001001111101100100011100111;
		b = 32'b10011100000001000100110110110001;
		correct = 32'b01011100101110001001010000111101;
		#400 //-0.00018194654 * -4.377555e-22 = 4.156351e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011100110111110011011101000111;
		b = 32'b01001011100011011000100111011101;
		correct = 32'b00010000110010011101110101100000;
		#400 //1.4771191e-21 * 18551738.0 = 7.9621603e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010111101010110111001101111000;
		b = 32'b00001100010010011011110000000101;
		correct = 32'b01001010110110011001001000001101;
		#400 //1.1079764e-24 * 1.5541057e-31 = 7129350.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100011001011111011001001110100;
		b = 32'b11111110100100101001101011100010;
		correct = 32'b00100100000110010110011001101110;
		#400 //-3.241039e+21 * -9.743574e+37 = 3.3263348e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010011010100001110111011101101;
		b = 32'b11001011100101101000111011111101;
		correct = 32'b01000111001100011010000011011010;
		#400 //-897361700000.0 * -19734010.0 = 45472.85
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101010001110110000100100010000;
		b = 32'b10001010000000001100010011101101;
		correct = 32'b11011111101110011110101100001000;
		#400 //1.661208e-13 * -6.2000134e-33 = -2.679362e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111000101101111000111101011001;
		b = 32'b01010010100010010101001110110100;
		correct = 32'b10100101101010110001011111001011;
		#400 //-8.7528206e-05 * 294907400000.0 = -2.9679894e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111001010110101101111011111001;
		b = 32'b11100110001000111001010101110101;
		correct = 32'b10010010101010110100001011000000;
		#400 //0.00020873164 * -1.9312568e+23 = -1.0808072e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000100001011001101000001100011;
		b = 32'b10011000001011110110100111100101;
		correct = 32'b00101011011111000011010011000001;
		#400 //-2.031419e-36 * -2.2671683e-24 = 8.9601595e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110010000110101100110001101001;
		b = 32'b00011011101001111000100000010010;
		correct = 32'b01010101111011001000101100000010;
		#400 //9.010457e-09 * 2.7715766e-22 = 32510222000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110111000010100101001100111101;
		b = 32'b11001101110100101100000000110001;
		correct = 32'b11101000101010000000011000110110;
		#400 //2.8055673e+33 * -441976350.0 = -6.347777e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101110100101100101010101000100;
		b = 32'b01001110011110000100010001010111;
		correct = 32'b00011111100110110000010000000010;
		#400 //6.8363565e-11 * 1041307100.0 = 6.5651684e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111000110000110011010011100010;
		b = 32'b00011100011011011101010111111011;
		correct = 32'b11011011110100100001110101110001;
		#400 //-9.308175e-05 * 7.8693285e-22 = -1.1828423e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110101100100101000111111100000;
		b = 32'b11011100011000111101010111111101;
		correct = 32'b10011000101001001010110111101100;
		#400 //1.0919721e-06 * -2.5652041e+17 = -4.2568623e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101011101011110100100100110100;
		b = 32'b00111001111011000110100000010011;
		correct = 32'b01110001001111011101000001001111;
		#400 //4.2381542e+26 * 0.0004509097 = 9.3991194e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011111110101100110100001101010;
		b = 32'b01001011111011010001010110010001;
		correct = 32'b00010011011001111000001110101111;
		#400 //9.0805264e-20 * 31075106.0 = 2.9221224e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111000010111110011010010111;
		b = 32'b00010110011010100011010111000100;
		correct = 32'b01110000000110001110101010100011;
		#400 //35814.59 * 1.8919335e-25 = 1.8930152e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100010111001011010000001010;
		b = 32'b00101000011011101101000010001000;
		correct = 32'b01011011011011001001010111011100;
		#400 //882.8131 * 1.3256872e-14 = 6.6592867e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000001010010111011101011110111;
		b = 32'b00111110100000001011110111010110;
		correct = 32'b01000010010010101000111010001110;
		#400 //12.733146 * 0.25144833 = 50.639214
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000000110001001000000111101111;
		b = 32'b10110010101011011110111111110010;
		correct = 32'b01001101100100001001110000000010;
		#400 //-6.140861 * -2.0248965e-08 = 303267900.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111100000110010010101110100011;
		b = 32'b01001100011101111001011001010010;
		correct = 32'b01101111000111100110000000000100;
		#400 //3.181226e+36 * 64903496.0 = 4.9014707e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110001010100001011110111001010;
		b = 32'b11001101111110101100101111111100;
		correct = 32'b11100010110101010001001001110001;
		#400 //1.0336372e+30 * -525959040.0 = -1.9652427e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011100111111010100011000100000;
		b = 32'b10110110001011001001010011000110;
		correct = 32'b00100110001110111101100100100101;
		#400 //-1.6760262e-21 * -2.5716595e-06 = 6.5172944e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111010010011101001000100001001;
		b = 32'b01001101010100001110010101101110;
		correct = 32'b00101100011111010010010100100000;
		#400 //0.0007879888 * 219043550.0 = 3.597407e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011001011011000000001000101001;
		b = 32'b00010101011110001101001100001111;
		correct = 32'b11000011011100101101000001111101;
		#400 //-1.220135e-23 * 5.0249697e-26 = -242.8144
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101110000010110001110111100011;
		b = 32'b10111000011110000001100010111101;
		correct = 32'b01110101000011111000110001100111;
		#400 //-1.0763637e+28 * -5.9150847e-05 = 1.8196927e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010010001101101101001011100000;
		b = 32'b10110110001110001000001000111111;
		correct = 32'b11011011011111011010100101111101;
		#400 //196305490000.0 * -2.749395e-06 = -7.1399523e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000001000000110101101110100111;
		b = 32'b00001001011000100110000010100000;
		correct = 32'b00110111000101001000101111111101;
		#400 //2.4126657e-38 * 2.7249193e-33 = 8.854081e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000000101010010111101100001001;
		b = 32'b10000110110010100001110011101011;
		correct = 32'b10111001010101101010101011010001;
		#400 //1.5564336e-38 * -7.6026446e-35 = -0.00020472264
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011111001101011110000111111110;
		b = 32'b11011000011000001100010111100101;
		correct = 32'b00000110010011110010011010110010;
		#400 //-3.8515177e-20 * -988562200000000.0 = 3.8960802e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000101000011010110100011110000;
		b = 32'b01001100001001100000000000011111;
		correct = 32'b00111000010110100001001111001011;
		#400 //2262.5586 * 43516028.0 = 5.1993684e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100100111111000001111111000001;
		b = 32'b10101101110101110010101101101000;
		correct = 32'b01110110100101011111101111000101;
		#400 //-3.720694e+22 * -2.4461946e-11 = 1.5210131e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011000111101101110010101011111;
		b = 32'b11101001110100111111010111010011;
		correct = 32'b00101110100101010001100011100100;
		#400 //-2171720000000000.0 * -3.2030527e+25 = 6.780157e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100011100001110001101111111011;
		b = 32'b01011011011011100111111001111111;
		correct = 32'b00000111100100010000011011001100;
		#400 //1.464858e-17 * 6.713013e+16 = 2.182117e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110110111101101100010110001;
		b = 32'b00111001010001100110111101010011;
		correct = 32'b01000101000011111011111100100100;
		#400 //0.43524697 * 0.00018924223 = 2299.9463
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011101101011011111010100011011;
		b = 32'b00100110110110110100001100011000;
		correct = 32'b00110110010010110001101010111101;
		#400 //4.604615e-21 * 1.5214363e-15 = 3.026492e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100011111001010001001010100111;
		b = 32'b10101100100110000110010100001000;
		correct = 32'b10110110110000000110011101100110;
		#400 //2.483613e-17 * -4.3313166e-12 = -5.734083e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011100010010100001111100110100;
		b = 32'b00101101100011110010100111110110;
		correct = 32'b00101110001101001011011010010001;
		#400 //6.6876523e-22 * 1.6275852e-11 = 4.1089413e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001010100101111110110110110010;
		b = 32'b00010010101001110111111110100000;
		correct = 32'b10110111011010000011010000000101;
		#400 //-1.4630182e-32 * 1.0570644e-27 = -1.3840389e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100101000111011111010110010000;
		b = 32'b10110101001001101000000100101011;
		correct = 32'b11101111011100101101110010010001;
		#400 //4.6621335e+22 * -6.2027783e-07 = -7.516202e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110011001001011010010011110101;
		b = 32'b10010110011101000100000001110011;
		correct = 32'b11011100001011011001110010010111;
		#400 //3.8567084e-08 * -1.97305e-25 = -1.9546937e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011011110101011001000001100011;
		b = 32'b11101100110111010100101001000101;
		correct = 32'b00101110011101110000111111100010;
		#400 //-1.2022585e+17 * -2.1401867e+27 = 5.6175405e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101001101000001010101000101000;
		b = 32'b01011100001101000011100111101010;
		correct = 32'b01001100111001000011011011001100;
		#400 //2.427896e+25 * 2.029167e+17 = 119649890.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101000101110000000101001111001;
		b = 32'b01011001110110000001101011101111;
		correct = 32'b00001110010110100000010000110001;
		#400 //2.0432645e-14 * 7603526000000000.0 = 2.6872593e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000110100110000001011010000000;
		b = 32'b01110011110101001101111010100000;
		correct = 32'b00010010001101101110011100101101;
		#400 //19467.25 * 3.373054e+31 = 5.771402e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111010111111000011101101101;
		b = 32'b01101011001000010000010001111001;
		correct = 32'b10001011101100011011000101110111;
		#400 //-1.3323367e-05 * 1.9465818e+26 = -6.844494e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110111011100100010110000001101;
		b = 32'b11000000000110010001111001111001;
		correct = 32'b11110110110010100111000110101000;
		#400 //4.9118332e+33 * -2.392485 = -2.0530258e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001101011011100001010111110000;
		b = 32'b00101001100000000001111000001001;
		correct = 32'b10100011011011011101111000011111;
		#400 //-7.336582e-31 * 5.689552e-14 = -1.2894832e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100000011101011111001100010100;
		b = 32'b11010111011010111000010110101010;
		correct = 32'b11001000100001011010101011000001;
		#400 //7.0890124e+19 * -258959320000000.0 = -273750.03
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001001111011010111011101101101;
		b = 32'b11111010000110111101100011111110;
		correct = 32'b00001111010000110000100011101010;
		#400 //-1945325.6 * -2.0230178e+35 = 9.615959e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001000101001111010010100011010;
		b = 32'b00010001010100010101011110001111;
		correct = 32'b11110110110011010000001001101110;
		#400 //-343336.8 * 1.6514174e-28 = -2.0790432e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100101011010011011000111111100;
		b = 32'b11000000001100110011011010100010;
		correct = 32'b00100100101001101110100110100110;
		#400 //-2.0269832e-16 * -2.8002095 = 7.238684e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100101001001011011101001011000;
		b = 32'b00001000101011101101101110011000;
		correct = 32'b01011011111100101010001000101000;
		#400 //1.4374604e-16 * 1.052387e-33 = 1.3659047e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111110110001000100111000001100;
		b = 32'b11111000101110111001101011110110;
		correct = 32'b01000101100001011110111110000001;
		#400 //-1.3046696e+38 * -3.0440703e+34 = 4285.938
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000010110100010111101111000010;
		b = 32'b00101110100010111001101000000001;
		correct = 32'b01010011110000000001001100000111;
		#400 //104.741714 * 6.348345e-11 = 1649905900000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101001100000001000011100101010;
		b = 32'b10101110100110111111000110011110;
		correct = 32'b10111010010100101111111001100100;
		#400 //5.707789e-14 * -7.091504e-11 = -0.00080487714
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001111001011101010010011100100;
		b = 32'b01001101000100000110001010100101;
		correct = 32'b01000001100110101101001100101101;
		#400 //2930041900.0 * 151398990.0 = 19.353113
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101110111110110101111111000011;
		b = 32'b10100111111001101110011011000000;
		correct = 32'b11000110100010110101100101011010;
		#400 //1.1431169e-10 * -6.4088004e-15 = -17836.676
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000111101110001001010000011101;
		b = 32'b01010101110000010100010110101011;
		correct = 32'b10110001011101000111110000100000;
		#400 //-94504.23 * 26563120000000.0 = -3.557723e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101101001100000100110110101110;
		b = 32'b11010101001010110000001110000101;
		correct = 32'b11010111100000111111010110001111;
		#400 //3.4102044e+27 * -11751975000000.0 = -290181380000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111001010100011000110110101001;
		b = 32'b00100101010110000000010100110100;
		correct = 32'b11010011011110000101011000001111;
		#400 //-0.00019984566 * 1.8736776e-16 = -1066595700000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111101000100111101111011101;
		b = 32'b00100111110110100101100000101100;
		correct = 32'b11001111001111101000000101110111;
		#400 //-1.9369583e-05 * 6.060275e-15 = -3196155600.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000011111011000010011101100111;
		b = 32'b00100010011101110100010000011101;
		correct = 32'b00100000111101000111111011001111;
		#400 //1.387988e-36 * 3.35108e-18 = 4.1419123e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010101111100101011101110000010;
		b = 32'b10110010000111000011011001100110;
		correct = 32'b01100011010001101110010011101000;
		#400 //-33360894000000.0 * -9.092764e-09 = 3.6689498e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101001011111110110001111001011;
		b = 32'b11001001101110011101101110010101;
		correct = 32'b01011111001011111110001011111100;
		#400 //-1.9296709e+25 * -1522546.6 = 1.2673969e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111101010111101111100011100111;
		b = 32'b01111001101101000111001000011101;
		correct = 32'b10000011000111100010101010011000;
		#400 //-0.05443659 * 1.1711599e+35 = -4.648092e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100101110110101011101100101001;
		b = 32'b00101001110110100111101111111101;
		correct = 32'b01111011100000000010010100000010;
		#400 //1.2911605e+23 * 9.702653e-14 = 1.3307292e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011000000101000110110101100111;
		b = 32'b11101010000001000010110010010000;
		correct = 32'b00101101100011111011110101110001;
		#400 //-652790400000000.0 * -3.994716e+25 = 1.6341347e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110100011110000001010101000100;
		b = 32'b01100101101011101101010111111101;
		correct = 32'b01001110001101011010000000011000;
		#400 //7.8620663e+31 * 1.0320489e+23 = 761792000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111011011111110001010101011110;
		b = 32'b11011101101010100110100000011001;
		correct = 32'b11011101001111111001101011000011;
		#400 //1.3244691e+36 * -1.5348865e+18 = -8.629101e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111111011000001001101100001111;
		b = 32'b01100011110101000100001010110000;
		correct = 32'b11011011000001110111000111001111;
		#400 //-2.9855218e+38 * 7.83103e+21 = -3.8124256e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001000110000010100011011110110;
		b = 32'b10011111110011010111011000011110;
		correct = 32'b11101000011100001101000110011011;
		#400 //395831.7 * -8.7016286e-20 = -4.548938e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110101011011110011100110100100;
		b = 32'b11001000001011000000001010000011;
		correct = 32'b01101100101100100000010010010011;
		#400 //-3.0325392e+32 * -176138.05 = 1.7216832e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011111010010001110111001010110;
		b = 32'b00000100011000100111001010000001;
		correct = 32'b01011010011000110010011101011000;
		#400 //4.2548794e-20 * 2.661875e-36 = 1.598452e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010101101111101011100010000000;
		b = 32'b00111110001100000000100100111011;
		correct = 32'b01010111000010101010110101110100;
		#400 //26212454000000.0 * 0.17191021 = 152477580000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001001101000001001000000110111;
		b = 32'b10110101011011101011101101010000;
		correct = 32'b00010011101011000010110101101110;
		#400 //-3.8654218e-33 * -8.8934485e-07 = 4.34637e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111111001100011100100110100000;
		b = 32'b10010001110000011111000011110011;
		correct = 32'b01101100111010101010110101101100;
		#400 //-0.6944828 * -3.0598527e-28 = 2.2696608e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010010100010000011100001111000;
		b = 32'b00111100100111001010110000101011;
		correct = 32'b11010101010111101001010011110111;
		#400 //-292531470000.0 * 0.019125065 = -15295711000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000010101011100010011101011110;
		b = 32'b10110111110001110100010101100111;
		correct = 32'b10001010010111111011101101110011;
		#400 //2.5589598e-37 * -2.3754967e-05 = -1.0772315e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010110110010010100110000001110;
		b = 32'b10100010000010010001101111010100;
		correct = 32'b00110100001110111110110010010001;
		#400 //-3.2521299e-25 * -1.8581694e-18 = 1.7501795e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011110111111110110001101101011;
		b = 32'b01010111010000101001001111111001;
		correct = 32'b10000111001010000000000011001011;
		#400 //-2.7040294e-20 * 213940800000000.0 = -1.2639148e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110010010111101100001100011001;
		b = 32'b10011011011111101101010101010100;
		correct = 32'b01010110010111111100100000101110;
		#400 //-1.2966461e-08 * -2.1079318e-22 = 61512715000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110100011110111101100000000101;
		b = 32'b01011101101000110111101100110001;
		correct = 32'b01010110010001010010111101001111;
		#400 //7.9812494e+31 * 1.4725079e+18 = 54201745000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101101001011011000110000100001;
		b = 32'b00101110100111100010010000111010;
		correct = 32'b00111110000011000111100000110011;
		#400 //9.865026e-12 * 7.191443e-11 = 0.13717727
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100001110001100110110000110011;
		b = 32'b01010010111110000000100010100011;
		correct = 32'b00001110010011001100101110100111;
		#400 //1.3445642e-18 * 532648400000.0 = 2.5242996e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001110001101011111111001011010;
		b = 32'b00101010010101000000000001100101;
		correct = 32'b11100011010110111100001110100011;
		#400 //-763336300.0 * 1.882952e-13 = -4.053934e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110110000101100000011011011110;
		b = 32'b11100000010110101110111100100110;
		correct = 32'b01010101001011110110110100110011;
		#400 //-7.607264e+32 * -6.310348e+19 = 12055221000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001111101111011111001000110001;
		b = 32'b00011110101011111010011011111011;
		correct = 32'b10110000100010100110101010000011;
		#400 //-1.8730128e-29 * 1.8597907e-20 = -1.0071094e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011010011010010101000001111110;
		b = 32'b01010010000110011011100100101000;
		correct = 32'b00000111110000100100010111010101;
		#400 //4.8248292e-23 * 165059100000.0 = 2.923092e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110111110101110111010111111111;
		b = 32'b01000000011100111000011010111111;
		correct = 32'b00110110111000100111111100111110;
		#400 //2.5684943e-05 * 3.8050992 = 6.750138e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101000101010000101010001000001;
		b = 32'b10111100011000010001010101111011;
		correct = 32'b00101011101111110111001100100010;
		#400 //-1.8688286e-14 * -0.0137380315 = 1.3603322e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101011001110100001011001011000;
		b = 32'b11100000001110010010001000010101;
		correct = 32'b11001010100000001010100011100010;
		#400 //2.2496572e+26 * -5.3360993e+19 = -4215921.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100010101011111110000001100101;
		b = 32'b00101001011010101001001111010110;
		correct = 32'b01111000101111111111000000110010;
		#400 //1.6221748e+21 * 5.2086665e-14 = 3.1143764e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011010000011100110101000001110;
		b = 32'b00111100010100001011010010001100;
		correct = 32'b11011101001011101010111111010010;
		#400 //-1.0021514e+16 * 0.012738358 = -7.867194e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011111111000001111010110011100;
		b = 32'b10100000101110011001001100000010;
		correct = 32'b11111110100110110010101001111100;
		#400 //3.2420068e+19 * -3.14375e-19 = -1.0312547e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011101111000001000110101010000;
		b = 32'b10110100011001110011110000001100;
		correct = 32'b10101000111110001001101000001011;
		#400 //5.943842e-21 * -2.1535396e-07 = -2.7600336e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100000011111010000110011011000;
		b = 32'b01001101001100101001010101101110;
		correct = 32'b10010010101101010101111110110111;
		#400 //-2.1434183e-19 * 187258600.0 = -1.1446301e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110101110101001110110001111100;
		b = 32'b10111000101001000111010010000100;
		correct = 32'b10111100101001011011100101110111;
		#400 //1.5864057e-06 * -7.841832e-05 = -0.020230038
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000100101100111110000000001001;
		b = 32'b00100011101100101000110100100110;
		correct = 32'b11100000100000001111001011110001;
		#400 //-1439.0011 * 1.9358577e-17 = -7.433403e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101110101110011011011100110101;
		b = 32'b10110111101101010101111111110100;
		correct = 32'b00110110100000110001000000111100;
		#400 //-8.44537e-11 * -2.1621563e-05 = 3.905994e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000001001111000001100111000000;
		b = 32'b00101110001000110010100111100011;
		correct = 32'b00010010100100111001000000010001;
		#400 //3.454862e-38 * 3.7099112e-11 = 9.312519e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010101010011101100100101101001;
		b = 32'b11111001000010000011011000010000;
		correct = 32'b00011011110000100101001000110011;
		#400 //-14210278000000.0 * -4.4203056e+34 = 3.2147728e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110011110110110011010011110010;
		b = 32'b11000000010110111010000111000010;
		correct = 32'b11110010111111111000000100101011;
		#400 //3.4734707e+31 * -3.431748 = -1.01215785e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111110110000000110001010010;
		b = 32'b10111001111011001100110101011010;
		correct = 32'b00111101011010011001000000111100;
		#400 //-2.5754944e-05 * -0.00045166427 = 0.05702232
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000000011101001110110000101011;
		b = 32'b10011001011000100011000100011100;
		correct = 32'b10100110100001000101010010110110;
		#400 //1.0737639e-38 * -1.1693844e-23 = -9.182301e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101111011111101101010111100100;
		b = 32'b00110100001011000101001011101110;
		correct = 32'b10111010101111010100100111011101;
		#400 //-2.3177155e-10 * 1.6048918e-07 = -0.0014441569
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110001000100011101110111010110;
		b = 32'b11100001111001010111001101110001;
		correct = 32'b11001110101000101011111010001011;
		#400 //7.2229615e+29 * -5.2907785e+20 = -1365198200.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010000010011000100000001100010;
		b = 32'b11010010111110111100010111110001;
		correct = 32'b00111100110011111010111000110100;
		#400 //-13707086000.0 * -540678850000.0 = 0.025351621
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010010111011110100001001011001;
		b = 32'b11000001011100111110001011001010;
		correct = 32'b01010000111110110010010010111010;
		#400 //-513805160000.0 * -15.242868 = 33707905000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011001110101100001110110100011;
		b = 32'b01000001001000001110110011111101;
		correct = 32'b10011000001010100100111010100111;
		#400 //-2.2139052e-23 * 10.057858 = -2.2011694e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101010000011000101101110011010;
		b = 32'b01001000111100100110111100001100;
		correct = 32'b00100000100101000011011001000111;
		#400 //1.2466279e-13 * 496504.38 = 2.5108093e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010101111010001101110110111011;
		b = 32'b10001101010000011000111000100101;
		correct = 32'b11001000000110011111111100100110;
		#400 //9.405388e-26 * -5.9643817e-31 = -157692.6
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111000010001100001011100100101;
		b = 32'b00000111100001100001011010111111;
		correct = 32'b01110000001111010001100001100110;
		#400 //4.7228434e-05 * 2.0175448e-34 = 2.3408865e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000000111001011001010111100000;
		b = 32'b00011011110000101110111110011011;
		correct = 32'b00100100100101101100000001110011;
		#400 //2.1084094e-38 * 3.224945e-22 = 6.537815e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000110111110000000001111111111;
		b = 32'b10000001011001111100110011001100;
		correct = 32'b01000101000010001111010001001011;
		#400 //-9.3293103e-35 * -4.2574934e-38 = 2191.2683
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101010100101101001110101010111;
		b = 32'b00010100000111110000000000110010;
		correct = 32'b11010101111100100111111101110010;
		#400 //-2.675453e-13 * 8.027487e-27 = -33328648000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101101100101110011010000011010;
		b = 32'b11000100001000010100110000001001;
		correct = 32'b01101000111011111111101011110011;
		#400 //-5.849403e+27 * -645.18805 = 9.066198e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100111110100110100111000010011;
		b = 32'b11101001100101010101010100110101;
		correct = 32'b10111101101101010001111010000001;
		#400 //1.9957191e+24 * -2.256654e+25 = -0.08843709
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101111101110111101010010100010;
		b = 32'b10010011101010011000010111010100;
		correct = 32'b01011011100011011101001011010011;
		#400 //-3.4166187e-10 * -4.2793562e-27 = 7.983955e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010010000011110010100100001010;
		b = 32'b11001010101101111111001111111100;
		correct = 32'b11000110110001110011101011111010;
		#400 //153717210000.0 * -6027774.0 = -25501.488
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001011110011110100111111001001;
		b = 32'b00110000001000010101100110100001;
		correct = 32'b01011011001001000111011000101001;
		#400 //27172754.0 * 5.869883e-10 = 4.6291815e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001000101101000000110101100101;
		b = 32'b10001100100010100110010010000111;
		correct = 32'b10111011101001101000011111111011;
		#400 //1.0836505e-33 * -2.132277e-31 = -0.005082128
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100101000010101001100001011010;
		b = 32'b11110011111101110010111011111101;
		correct = 32'b10110000100011111000100111011010;
		#400 //4.090606e+22 * -3.9167797e+31 = -1.0443799e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110100010010010111011010011101;
		b = 32'b01011100010100010010111110111000;
		correct = 32'b10010111011101101000110001110001;
		#400 //-1.8762735e-07 * 2.3552295e+17 = -7.966415e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101110001011011000011100111000;
		b = 32'b11000110001000011111100010111100;
		correct = 32'b10100111100010010010000111111010;
		#400 //3.9455744e-11 * -10366.184 = -3.8061976e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010101010001100110010101100101;
		b = 32'b10111110001010010111011000100000;
		correct = 32'b00010110100101011101101011110111;
		#400 //-4.0065768e-26 * -0.16548967 = 2.4210435e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101110101100111001000100110100;
		b = 32'b11011100011011111001000111110100;
		correct = 32'b11010001101111111110000111001101;
		#400 //2.7786678e+28 * -2.6973199e+17 = -103015880000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001110001111110100010000001111;
		b = 32'b01010110010111001011011010000000;
		correct = 32'b10110111010111011101100001010100;
		#400 //-802227140.0 * 60669097000000.0 = -1.3222994e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100100010001111111100010011000;
		b = 32'b11000000011111110010001111010111;
		correct = 32'b10100011010010001010010100100110;
		#400 //4.3361814e-17 * -3.9865625 = -1.0876993e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001111111001110111111000111011;
		b = 32'b01101000100011100001010001000111;
		correct = 32'b10100110110100001000110110110010;
		#400 //-7767619000.0 * 5.367601e+24 = -1.4471306e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001011110011110101110000110111;
		b = 32'b00101101110000010001100111011101;
		correct = 32'b00011101100010010111001110110001;
		#400 //7.987225e-32 * 2.1953045e-11 = 3.638322e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101101011100100000110100010001;
		b = 32'b00111000101100000001000100000110;
		correct = 32'b11110100001011111111100001111011;
		#400 //-4.681948e+27 * 8.395505e-05 = -5.576732e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000100011100101000000010001111;
		b = 32'b00000101001100001100011101111110;
		correct = 32'b10111110101011111001011001111001;
		#400 //-2.8505995e-36 * 8.312121e-36 = -0.3429449
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010001011011110110101000000110;
		b = 32'b00111110110101100011111011111011;
		correct = 32'b01010010000011110000100101011100;
		#400 //64267248000.0 * 0.41844925 = 153584340000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011001001010100110001101101010;
		b = 32'b01000000000101001001000100111111;
		correct = 32'b01011000100100101100110011010101;
		#400 //2997503300000000.0 * 2.321365 = 1291267600000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011110010101011010010101011100;
		b = 32'b00111110010101010101101000101111;
		correct = 32'b11011111100000000010110100011010;
		#400 //-3.848703e+18 * 0.20835184 = -1.8472134e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110011110100011011100101111011;
		b = 32'b10000001001011101101000100001001;
		correct = 32'b11110010000110011000111100111011;
		#400 //9.7660596e-08 * -3.2108728e-38 = -3.041559e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100100101111010001000100100101;
		b = 32'b00110110001001111010010000101000;
		correct = 32'b00101110000100000101101111111011;
		#400 //8.199473e-17 * 2.498049e-06 = 3.2823504e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110110000110001101000010111101;
		b = 32'b01110101000000110100101110001101;
		correct = 32'b01000000100101001111101011101100;
		#400 //7.7486605e+32 * 1.6643634e+32 = 4.65563
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100010010000101100111100111001;
		b = 32'b11100001011010100111010101000010;
		correct = 32'b11000000010101001011010101100010;
		#400 //8.984001e+20 * -2.7031171e+20 = -3.3235707
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110000101110010011011111000;
		b = 32'b00110110100110001010010110110110;
		correct = 32'b01000110111111010111111000011101;
		#400 //0.14760959 * 4.5492443e-06 = 32447.057
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111001111111001110111001101001;
		b = 32'b10110111101101010000010000010010;
		correct = 32'b01000001101100101101101001010011;
		#400 //-0.00048242815 * -2.1578777e-05 = 22.356604
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111001010111011001111100111111;
		b = 32'b11100101111111101000010011000001;
		correct = 32'b10010010110111101110100101111010;
		#400 //0.00021135526 * -1.5024125e+23 = -1.4067726e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000001000010111101010011101111;
		b = 32'b01101001101110000000001001001001;
		correct = 32'b10010110110000101000101000000011;
		#400 //-8.739486 * 2.7806643e+25 = -3.1429488e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100110001010110111110110000111;
		b = 32'b11010100100101101000000110110010;
		correct = 32'b10010001000100011101100010001000;
		#400 //5.9497664e-16 * -5171368000000.0 = -1.1505207e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111001001000011111111001110001;
		b = 32'b00010111001111010101111110101001;
		correct = 32'b11100001010110101111110011000100;
		#400 //-0.00015448943 * 6.1189934e-25 = -2.5247524e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001010101000000011111001101000;
		b = 32'b00011111001001110001111000001110;
		correct = 32'b00101010111101010111100001111000;
		#400 //1.5430914e-32 * 3.5388486e-20 = 4.3604335e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100001011110111011111110100011;
		b = 32'b00110100110100001010100100010001;
		correct = 32'b00101100000110100110111010001111;
		#400 //8.5295737e-19 * 3.886603e-07 = 2.1946089e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100111000110101100111010001011;
		b = 32'b00101001001001010001111001000101;
		correct = 32'b10111101011100000000001101011011;
		#400 //-2.148376e-15 * 3.6663614e-14 = -0.05859695
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111000101001000111110110000010;
		b = 32'b01100011010110110010110110111100;
		correct = 32'b10010100110000000001111111000111;
		#400 //-7.843507e-05 * 4.0431325e+21 = -1.939958e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111111110010011011100100010010;
		b = 32'b01010100000001000111100110100101;
		correct = 32'b11111111110010011011100100010010;
		#400 //nan * 2275906200000.0 = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100111010011101100111101011101;
		b = 32'b11111101011111010011110101110101;
		correct = 32'b00101001010100010001000001011110;
		#400 //-9.766327e+23 * -2.1038362e+37 = 4.642152e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001010001001000101011110110001;
		b = 32'b10001010110011001001001111001111;
		correct = 32'b10111110110011011010011011011000;
		#400 //7.912806e-33 * -1.9700085e-32 = -0.40166354
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101110000001001001100110001100;
		b = 32'b01000001110100101011001111001001;
		correct = 32'b01101011101000010001101101010000;
		#400 //1.0259412e+28 * 26.337786 = 3.8953207e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110001000011100001000001111111;
		b = 32'b01000010101011101001001011010001;
		correct = 32'b10101101110100000101001111100100;
		#400 //-2.0673097e-09 * 87.28675 = -2.3684117e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101111000011100111111001100101;
		b = 32'b01111001000110010100000101000010;
		correct = 32'b10110101011011100000011000111001;
		#400 //-4.4099673e+28 * 4.9734063e+34 = -8.8670964e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101110101111100111111111110110;
		b = 32'b01011010010001010111000110101110;
		correct = 32'b10010011111101101111111100010000;
		#400 //-8.66293e-11 * 1.3893891e+16 = -6.235064e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001001100000100111101001010000;
		b = 32'b01000000111001011010011101100011;
		correct = 32'b11001000000100010111001001000011;
		#400 //-1068874.0 * 7.176683 = -148937.05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101100001010111100010001010100;
		b = 32'b00101010010000001100001111100001;
		correct = 32'b01000001011001000001110100001101;
		#400 //2.4409546e-12 * 1.7120985e-13 = 14.257092
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101011100111011110001000110001;
		b = 32'b00111100111010000010110010101011;
		correct = 32'b00101110001011100001010111011110;
		#400 //1.1218302e-12 * 0.028341612 = 3.958244e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001111100011011110010111101110;
		b = 32'b00110001010110110111010100111101;
		correct = 32'b01011101101001011000011010010011;
		#400 //4761312000.0 * 3.1935337e-09 = 1.4909228e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000011100010101111101100101100;
		b = 32'b00001111111011100101000001100000;
		correct = 32'b10110011000101010100101110011101;
		#400 //-8.168577e-37 * 2.3499571e-29 = -3.4760536e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001101111011110111100010101101;
		b = 32'b11101101000001011111101101010111;
		correct = 32'b00100000011001001100011110100110;
		#400 //-502207900.0 * -2.5915848e+27 = 1.9378409e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001110010010011000100111101011;
		b = 32'b00011010110010110011101101110001;
		correct = 32'b00110010111111011101110111101010;
		#400 //2.4841568e-30 * 8.4054865e-23 = 2.9553991e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101011011101101001110011010011;
		b = 32'b00111000000101111011111111011111;
		correct = 32'b01110010110100000000010000111111;
		#400 //2.9813633e+26 * 3.61799e-05 = 8.240386e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010000001001101110011101101101;
		b = 32'b11100011110001100000100011010010;
		correct = 32'b10101011110101111100000111101110;
		#400 //11200738000.0 * -7.306182e+21 = -1.5330495e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010011110110111100010000011010;
		b = 32'b11011010011011011000011001001010;
		correct = 32'b10111000111011001101110000110010;
		#400 //1887775800000.0 * -1.6714305e+16 = -0.000112943715
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010000100111111110010000011110;
		b = 32'b11001010110100011000110111010101;
		correct = 32'b00000101010000110101010001100100;
		#400 //-6.306591e-29 * -6866666.5 = 9.184356e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110110010010110100100101101101;
		b = 32'b00111001111111000101100001100110;
		correct = 32'b01111011110011100011101100100011;
		#400 //1.0307866e+33 * 0.00048131048 = 2.1416252e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111001111100000101101110000000;
		b = 32'b00010110110011101001001010101101;
		correct = 32'b11100010100101001110111100011111;
		#400 //-0.0004584454 * 3.337366e-25 = -1.3736743e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011110010101001111010011010101;
		b = 32'b01100001101011111110111000101100;
		correct = 32'b10111100000110101111000001001101;
		#400 //-3.836281e+18 * 4.056678e+20 = -0.009456706
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001100101011010010101011001010;
		b = 32'b00011011110010101010001001000111;
		correct = 32'b10110000010110101100010111011000;
		#400 //-2.6680623e-31 * 3.3522966e-22 = -7.958909e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101101011011110010000101110011;
		b = 32'b11010101111110000001101011100100;
		correct = 32'b10010110111101101011110101110100;
		#400 //1.3593004e-11 * -34099297000000.0 = -3.9863005e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010000000000110011101010111000;
		b = 32'b11100010110100010001100010001010;
		correct = 32'b10101100101000001010101010100110;
		#400 //8806654000.0 * -1.9285689e+21 = -4.5664193e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001011011111110110000100000010;
		b = 32'b00011001000010011011011111100000;
		correct = 32'b00110001111011010101101110011001;
		#400 //4.9184194e-32 * 7.119867e-24 = 6.9080213e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000000111011100000110010101110;
		b = 32'b01111011100110000111111011010000;
		correct = 32'b10000100110001111100111111000100;
		#400 //-7.439048 * 1.5836024e+36 = -4.6975478e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111101001100100010000001000101;
		b = 32'b01111011001011110100010101011101;
		correct = 32'b10000001100000100001010111000111;
		#400 //-0.043487806 * 9.100588e+35 = -4.7785707e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111000011100000001010110011010;
		b = 32'b00101011000011101110000001101010;
		correct = 32'b01001100110101110001011000010111;
		#400 //5.7240577e-05 * 5.075997e-13 = 112767160.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100010100000111010011000100100;
		b = 32'b11100000011010111000000111011001;
		correct = 32'b10000001100011110001101011000000;
		#400 //3.568353e-18 * -6.7880334e+19 = -5.256829e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011010110011100011100001111100;
		b = 32'b11000101100110001011001110100111;
		correct = 32'b11010100101011001101110010000101;
		#400 //2.9022975e+16 * -4886.4565 = -5939472600000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010111001100001000001101001100;
		b = 32'b11000001101011010011011001101100;
		correct = 32'b10010101000000100111000001011000;
		#400 //5.7034387e-25 * -21.651573 = -2.6341915e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000011011001010000011000111101;
		b = 32'b01110001110001000100101111011110;
		correct = 32'b10010001000101010101011101010100;
		#400 //-229.02437 * 1.944025e+30 = -1.1780938e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110101000011110110101100111000;
		b = 32'b01100011010001000000000001010100;
		correct = 32'b10010001001110110101001001000010;
		#400 //-5.3427675e-07 * 3.6155855e+21 = -1.4777047e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000010000001111101100101000101;
		b = 32'b00000111100000001010011010100010;
		correct = 32'b01111010000001110010100101010000;
		#400 //33.962177 * 1.9357237e-34 = 1.754495e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101000100010001100001111000000;
		b = 32'b11000110001001101100100100111111;
		correct = 32'b10100001110100011110101110001000;
		#400 //1.5183926e-14 * -10674.312 = -1.4224735e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001100100001001000110011001001;
		b = 32'b11000000001110011000011100100111;
		correct = 32'b01001011101101101110011000000101;
		#400 //-69494344.0 * -2.898874 = 23972874.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101000000111011001101100001010;
		b = 32'b01011011101010010100110010010110;
		correct = 32'b11001011111011100101000101101001;
		#400 //-2.977086e+24 * 9.530696e+16 = -31236818.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111001110110000100011100110110;
		b = 32'b11101110011001100010110001111100;
		correct = 32'b01001010111100001000101110010111;
		#400 //-1.4037256e+35 * -1.7808833e+28 = 7882187.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100110010010011110110110110111;
		b = 32'b11011001101110010101001111011111;
		correct = 32'b10001100000010110111011100111100;
		#400 //7.005805e-16 * -6520636000000000.0 = -1.0744051e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110111000110110001100101011010;
		b = 32'b01110101110101001000101101001101;
		correct = 32'b00000000101110101100111101010110;
		#400 //9.244623e-06 * 5.3886342e+32 = 1.715578e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100111010110110111100010000111;
		b = 32'b00110101101101100100010001111111;
		correct = 32'b11110001000110100010000001100011;
		#400 //-1.0364216e+24 * 1.3579992e-06 = -7.631975e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000011011010111111110111101001;
		b = 32'b00111011100110111010011111001010;
		correct = 32'b00000111010000100001000000011111;
		#400 //6.9351768e-37 * 0.0047502266 = 1.4599675e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010111100111101110101110100010;
		b = 32'b01110100110010110110001011100101;
		correct = 32'b00100010010010000000100000000101;
		#400 //349469740000000.0 * 1.2891139e+32 = 2.71093e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000010111000111111000111011011;
		b = 32'b10111100000000001010011100101101;
		correct = 32'b10000110011000101100100110101000;
		#400 //3.349347e-37 * -0.007852358 = -4.265403e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010000100010000010111100010100;
		b = 32'b10011101111100110000110000111000;
		correct = 32'b10110010000011110111000011111000;
		#400 //5.3715077e-29 * -6.43342e-21 = -8.349382e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000100010000010011111101101100;
		b = 32'b11110101010011101100010111011011;
		correct = 32'b00001110011011110100000101000001;
		#400 //-772.99097 * -2.6211576e+32 = 2.9490443e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110111111101010100000010011101;
		b = 32'b11111000101000100011100101001110;
		correct = 32'b10111110110000011000001100100101;
		#400 //9.948619e+33 * -2.6322324e+34 = -0.37795368
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010010110011010010111011101001;
		b = 32'b01101001101100001110100101000100;
		correct = 32'b10101000100101000111010010100001;
		#400 //-440627660000.0 * 2.6734064e+25 = -1.648188e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110111010110010111111001110110;
		b = 32'b11000111100010100100000101110010;
		correct = 32'b11101111010010010101110001001100;
		#400 //4.411302e+33 * -70786.89 = -6.2318067e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110100011111100011100111000;
		b = 32'b01001011110101111010000110101101;
		correct = 32'b10101010001010101011000111101001;
		#400 //-4.284924e-06 * 28263258.0 = -1.5160758e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010010010111100101010010111011;
		b = 32'b11100001101100111010010101101111;
		correct = 32'b00110000000111100110100111010011;
		#400 //-238726070000.0 * -4.14236e+20 = 5.763045e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111111110011100111101001001;
		b = 32'b00110010001011001100110000001101;
		correct = 32'b01010101001110010000110000100000;
		#400 //127902.57 * 1.00581135e-08 = 12716358000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011110110110000000011110011001;
		b = 32'b00010101001101100100010001111010;
		correct = 32'b01001001000101111011010111000010;
		#400 //2.2873032e-20 * 3.6808626e-26 = 621404.1
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001111010000111000010101111110;
		b = 32'b00011010111011111011000110110001;
		correct = 32'b00110011110100001101001010000111;
		#400 //9.639952e-30 * 9.913516e-23 = 9.7240495e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111110100010101001100011100011;
		b = 32'b11010001010000110010000010000101;
		correct = 32'b00101100101101011101010110110110;
		#400 //-0.27069768 * -52379013000.0 = 5.168056e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001010100001101101100011000000;
		b = 32'b01011010010010000000010101010001;
		correct = 32'b00101111101011001001010111111001;
		#400 //4418656.0 * 1.407521e+16 = 3.139318e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000001101100110000010111100101;
		b = 32'b01110000100000101110010110000100;
		correct = 32'b00010000101011110000111110111111;
		#400 //22.377878 * 3.2408415e+29 = 6.904959e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001100100111010000111001110100;
		b = 32'b01100001001011010110111001100011;
		correct = 32'b10101010111001111101010001010101;
		#400 //-82342820.0 * 1.9995256e+20 = -4.1181178e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011011001101111101100111001010;
		b = 32'b01001101010110001010101011001100;
		correct = 32'b01001101010110010011100111101001;
		#400 //5.1749382e+16 * 227192000.0 = 227778190.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001111111110010100000101011110;
		b = 32'b00010100000111100001001110100011;
		correct = 32'b01111011010010011101010010010101;
		#400 //8363621400.0 * 7.980834e-27 = 1.04796334e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000001110000100010100010011101;
		b = 32'b10010100100110000100111110001001;
		correct = 32'b10101100101000110010101100100011;
		#400 //7.132262e-38 * -1.5379449e-26 = -4.6375278e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011100001010001101010010101101;
		b = 32'b01000101111110000001001001001100;
		correct = 32'b10010101101011100011101000001001;
		#400 //-5.5861414e-22 * 7938.287 = -7.0369604e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000100100011011101011101011111;
		b = 32'b00110101111111111101011001101010;
		correct = 32'b11001110000011011110111001101101;
		#400 //-1134.7303 * 1.9061383e-06 = -595303230.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001001111101110111000010100110;
		b = 32'b01101011010010101110100010101101;
		correct = 32'b10011110000111000001011101100011;
		#400 //-2027028.8 * 2.453018e+26 = -8.2634075e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100001011000110111101010000001;
		b = 32'b00011011100100101011100010101101;
		correct = 32'b11000101010001100111001111100010;
		#400 //-7.7072724e-19 * 2.4273018e-22 = -3175.2427
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010101000110100001000101000001;
		b = 32'b11100010101101101011011011011110;
		correct = 32'b10110001110101111101110011101011;
		#400 //10587431000000.0 * -1.6852422e+21 = -6.282439e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101000111101101110100010111010;
		b = 32'b10110010100010110010110010010111;
		correct = 32'b00110101111000110001010111000000;
		#400 //-2.7412415e-14 * -1.6202007e-08 = 1.6919148e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001110110110001011000010111100;
		b = 32'b11000110111000100011011100110111;
		correct = 32'b10000111011101010011100001110110;
		#400 //5.34183e-30 * -28955.607 = -1.8448344e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110101111101010110110011101110;
		b = 32'b10101000111010100001010101010010;
		correct = 32'b11001100100001100011001110111100;
		#400 //1.8285625e-06 * -2.5988465e-14 = -70360540.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000111001110100000011010001111;
		b = 32'b00101011000010001111110000001111;
		correct = 32'b00011011101011011101001100010010;
		#400 //1.3995012e-34 * 4.866671e-13 = 2.875685e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100111010101101001101001111110;
		b = 32'b00010011011101000100101011010110;
		correct = 32'b11010011011000001110001101101001;
		#400 //-2.9782216e-15 * 3.0834027e-27 = -965888000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110101100110010001110111000001;
		b = 32'b10100110100011111010101001000110;
		correct = 32'b01001110100010000110101110101010;
		#400 //-1.1408048e-06 * -9.968771e-16 = 1144378600.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101000001101100101111110011010;
		b = 32'b10011001010110100010000100111110;
		correct = 32'b11001110010101100000100100101011;
		#400 //1.012376e-14 * -1.1277049e-23 = -897731260.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101111101101111001101001001111;
		b = 32'b00111110000001100111000110100110;
		correct = 32'b01110001001011101100110101111001;
		#400 //1.1364461e+29 * 0.13129291 = 8.655807e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010011011100110110110111101101;
		b = 32'b10010111010001100000111010111010;
		correct = 32'b11111011100111010101001010100010;
		#400 //1045521300000.0 * -6.399584e-25 = -1.6337332e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100101000111110110011101110000;
		b = 32'b00011001100001010011100011101100;
		correct = 32'b11001011000110010010011111000110;
		#400 //-1.3826098e-16 * 1.3774868e-23 = -10037190.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010011010100101100111101000001;
		b = 32'b11100101111011101111010010010100;
		correct = 32'b10101100111000011101100010111001;
		#400 //905420300000.0 * -1.4105436e+23 = -6.4189457e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001100100101010101101001100000;
		b = 32'b00011011101110011010111000111011;
		correct = 32'b00110000010011011110101000101110;
		#400 //2.3011477e-31 * 3.0718276e-22 = 7.4911355e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011100011001100010110000000011;
		b = 32'b01000100111111001010010110111000;
		correct = 32'b01010110111010010011100111110001;
		#400 //2.5915054e+17 * 2021.1787 = 128217530000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000010110110011000011011010100;
		b = 32'b11000001010100101110111001000101;
		correct = 32'b01000001000001000000000010101101;
		#400 //-108.763336 * -13.183171 = 8.250165
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111110010000101111110011110001;
		b = 32'b11101110011000000111101110101010;
		correct = 32'b00001111010111100101110100101100;
		#400 //-0.19041802 * -1.7368536e+28 = 1.0963389e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010001111111110011100100011010;
		b = 32'b01001110111000110000011001100111;
		correct = 32'b10000010100011111110011000000010;
		#400 //-4.0267098e-28 * 1904423800.0 = -2.114398e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000100110101101011000111100000;
		b = 32'b00111010000000100111101100001100;
		correct = 32'b11001010010100101001110011110110;
		#400 //-1717.5586 * 0.0004977442 = -3450685.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101011001110000110010111000101;
		b = 32'b01001111000010010100010011100100;
		correct = 32'b00011011101010111111001000110011;
		#400 //6.5511165e-13 * 2302993400.0 = 2.8446095e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000000010100000111010100011001;
		b = 32'b11110101110100011010100110111111;
		correct = 32'b10001001111111101000011100100011;
		#400 //3.257147 * -5.3155903e+32 = -6.1275358e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000010111001101001101000100001;
		b = 32'b10111101011100111000011111011101;
		correct = 32'b11000100111100100110100011001101;
		#400 //115.30103 * -0.05945574 = -1939.275
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011010000001111000110101111010;
		b = 32'b00110000100110100101110100110001;
		correct = 32'b00101000111000001100110110001001;
		#400 //2.803163e-23 * 1.1231461e-09 = 2.4958132e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010101100011110101101001110001;
		b = 32'b11000001101101100000100010010100;
		correct = 32'b00010011010010011001101001001001;
		#400 //-5.789993e-26 * -22.754189 = 2.5445835e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001011011100111011010010010011;
		b = 32'b00111101010011011111001001101000;
		correct = 32'b00001101100101110111011110110110;
		#400 //4.6935947e-32 * 0.050280005 = 9.334913e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000010110100101011101010010101;
		b = 32'b10110011000010010001111110110011;
		correct = 32'b01001111010001001011010100100010;
		#400 //-105.36442 * -3.192663e-08 = 3300205000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001000001100010011010100000000;
		b = 32'b00011111100010011001110100111011;
		correct = 32'b00101000001001001101001110100111;
		#400 //5.33263e-34 * 5.828187e-20 = 9.149724e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011111110000010000101000011101;
		b = 32'b10000101010001101111011101000110;
		correct = 32'b01011001111110000101111111110001;
		#400 //-8.175541e-20 * -9.355332e-36 = 8738910400000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101000010010101100001100000001;
		b = 32'b01010001100101101101010110100110;
		correct = 32'b00010110001011000001000011100110;
		#400 //1.1255537e-14 * 80978690000.0 = 1.3899382e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111011100001100110000011011010;
		b = 32'b01110100111100000101011010001110;
		correct = 32'b11000110000011110010001010011111;
		#400 //-1.3954643e+36 * 1.5233237e+32 = -9160.655
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000100110111110111101001100111;
		b = 32'b10101101110010101111001110110110;
		correct = 32'b01010110100011001111001000010110;
		#400 //-1787.8251 * -2.307297e-11 = 77485690000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110111110001110111111010000000;
		b = 32'b11011001101101001000100101011011;
		correct = 32'b10011101100011010111000011011110;
		#400 //2.3781555e-05 * -6352065000000000.0 = -3.743909e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011111011000111010001110010011;
		b = 32'b11101001010101010000100111111001;
		correct = 32'b10110101100010001100010110101001;
		#400 //1.6403116e+19 * -1.6096768e+25 = -1.0190316e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001110101100010011111100000101;
		b = 32'b10110010000111010000101010101100;
		correct = 32'b10011100000100000111011111010100;
		#400 //4.3694554e-30 * -9.141029e-09 = -4.780048e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011101111000110011101010111101;
		b = 32'b01010100111110011011100111111101;
		correct = 32'b10001000011010001111000000010010;
		#400 //-6.0147134e-21 * 8580538000000.0 = -7.009716e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011110000101100011111101000011;
		b = 32'b01010111101101010011101100000101;
		correct = 32'b00000101110101000011101111100000;
		#400 //7.954016e-21 * 398530180000000.0 = 1.9958379e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001010010010011111001010011011;
		b = 32'b10101111100100100000001101110000;
		correct = 32'b11011010001100010000100010100011;
		#400 //3308710.8 * -2.6559688e-10 = -1.2457642e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010111100110001011010000101100;
		b = 32'b00101011110101101111101111111101;
		correct = 32'b10101011001101011101011001011010;
		#400 //-9.868252e-25 * 1.5275555e-12 = -6.460159e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011001101000100011111011010011;
		b = 32'b01011110010010101001111010101000;
		correct = 32'b00111010110011001111110100110000;
		#400 //5708503000000000.0 * 3.650073e+18 = 0.0015639421
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000101000001111000101010000011;
		b = 32'b10001100110111000100000111001001;
		correct = 32'b11110111100111011000100101011000;
		#400 //2168.657 * -3.393596e-31 = -6.3904396e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110000000011100100100111011111;
		b = 32'b10101010010101111100011100101010;
		correct = 32'b11000101001010001100111111010010;
		#400 //5.1764276e-10 * -1.9164935e-13 = -2700.9888
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100101110100010100101001111101;
		b = 32'b10110011101100011100000101110101;
		correct = 32'b11110001100101101011010101001110;
		#400 //1.2354358e+23 * -8.2773944e-08 = -1.492542e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011110011110111100000000011111;
		b = 32'b11010000000010101110010111110000;
		correct = 32'b00001101111001111111111101101001;
		#400 //-1.3327559e-20 * -9321300000.0 = 1.4297962e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101101001101011011111000111011;
		b = 32'b01011110001111100011000111111000;
		correct = 32'b11001110011101001001111110100100;
		#400 //-3.5154226e+27 * 3.426252e+18 = -1026025700.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110000111110101111100000000010;
		b = 32'b10001010100111101010111111100101;
		correct = 32'b11100101110010100110111110101000;
		#400 //1.8260382e-09 * -1.528101e-32 = -1.19497215e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110010101100101011111100010100;
		b = 32'b11011101011001100010101100000101;
		correct = 32'b00010100110001101100111010101001;
		#400 //-2.080882e-08 * -1.0365847e+18 = 2.0074404e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000100011001011111111101110001;
		b = 32'b00001110110111010101100110110100;
		correct = 32'b10110101000001010000000000100011;
		#400 //-2.7036114e-36 * 5.4567087e-30 = -4.954656e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111111000000001010110011110010;
		b = 32'b11000000001111000110100001000000;
		correct = 32'b11111110001011101101011011001110;
		#400 //1.7103917e+38 * -2.943863 = -5.810025e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001001110001101000101011000010;
		b = 32'b00110000001000111010100011001010;
		correct = 32'b00011001000110110100100000111101;
		#400 //4.7797253e-33 * 5.953892e-10 = 8.0279006e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010000101101100101001011110011;
		b = 32'b00111111101000110001100110101001;
		correct = 32'b10010000100011110001011000110010;
		#400 //-7.1914146e-29 * 1.2742206 = -5.643775e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110111010100011000100000000111;
		b = 32'b11100001110010011100101111000001;
		correct = 32'b11010101000001001110100000011001;
		#400 //4.2498008e+33 * -4.653097e+20 = -9133274000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001011101111000101000100001000;
		b = 32'b00001101001111111110001110011010;
		correct = 32'b00111101111110110011101111011110;
		#400 //7.253689e-32 * 5.9130385e-31 = 0.12267278
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011110110010000111111011100001;
		b = 32'b11000010111001010000001110010110;
		correct = 32'b01011011011000000001111100000011;
		#400 //-7.223616e+18 * -114.507 = 6.3084493e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111010011011011101110101111001;
		b = 32'b01001100010111011011010111101110;
		correct = 32'b01101101100010010101001110010010;
		#400 //3.0876659e+35 * 58120120.0 = 5.3125596e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111001100100101101000111010110;
		b = 32'b01011111111010010111110100010101;
		correct = 32'b11011001001000001111100110011100;
		#400 //-9.5291415e+34 * 3.3649254e+19 = -2831902800000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111111011001010110000100001101;
		b = 32'b10101101110010000011000001011000;
		correct = 32'b01010001000100101010101000000101;
		#400 //-0.8960121 * -2.2758836e-11 = 39369855000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011010011001010011011111101000;
		b = 32'b11011110010000000011100010101110;
		correct = 32'b10111011100110001010001011100001;
		#400 //1.612981e+16 * -3.462753e+18 = -0.0046580886
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100101011010010011011011010001;
		b = 32'b10101000110110101101101101001010;
		correct = 32'b00111100000010000110010110101001;
		#400 //-2.0228101e-16 * -2.4297963e-14 = 0.008325019
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000101100010011011000001100110;
		b = 32'b00001011100100101110001101100100;
		correct = 32'b11111001011011111111011110101011;
		#400 //-4406.05 * 5.6579294e-32 = -7.787389e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011010001001110111110110000100;
		b = 32'b01000010111011000101101110111001;
		correct = 32'b11010110101101010110100010110011;
		#400 //-1.1786082e+16 * 118.179146 = -99730640000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000100110101111111100111101100;
		b = 32'b10011100111011001000000111000101;
		correct = 32'b10100111011010011100011011110110;
		#400 //5.0775774e-36 * -1.5650715e-21 = -3.2443103e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111011010110101111111100111110;
		b = 32'b11101110110010101101101001101010;
		correct = 32'b11001100000010100010111111001111;
		#400 //1.13709764e+36 * -3.139001e+28 = -36224828.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110000010110111000010010000110;
		b = 32'b00001101001110011101011111110001;
		correct = 32'b01100010100101110011000101110000;
		#400 //7.9860063e-10 * 5.7267456e-31 = 1.3945104e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110010111110111101110001111110;
		b = 32'b01100110010101110001001100101000;
		correct = 32'b10001100000101011110010010100110;
		#400 //-2.9320514e-08 * 2.5391554e+23 = -1.1547349e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011001100011010010111001011111;
		b = 32'b01010110101101011111110111110111;
		correct = 32'b10000010010001101001011111010111;
		#400 //-1.4597787e-23 * 100051190000000.0 = -1.4590318e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100100100101110000011000110100;
		b = 32'b00110011101110001110010110001100;
		correct = 32'b01110000010100010001101000000111;
		#400 //2.2287243e+22 * 8.609922e-08 = 2.5885533e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110011111101101010010011000101;
		b = 32'b01101101000011011101000101011101;
		correct = 32'b11000110010111101001110010111100;
		#400 //-3.9082243e+31 * 2.7431557e+27 = -14247.184
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111000110011101100111101000100;
		b = 32'b10010000010011100010101110000110;
		correct = 32'b11101000000000000110010110101001;
		#400 //9.861452e-05 * -4.0659866e-29 = -2.4253528e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001010110010101101010100010001;
		b = 32'b11000000100101110101111000110100;
		correct = 32'b11001001101010111000010011110010;
		#400 //6646408.5 * -4.7302494 = -1405086.2
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000101010110001010111010101;
		b = 32'b11010001011001000000110110000010;
		correct = 32'b00011110110000000000110100100011;
		#400 //-1.2448093e-09 * -61217448000.0 = 2.0334224e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011110001011011000101101100000;
		b = 32'b00101111000011110101001110000000;
		correct = 32'b01101110100110101111110010101001;
		#400 //3.1262986e+18 * 1.303544e-10 = 2.398307e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101010010001010110110101001101;
		b = 32'b00010110001101110110000001011010;
		correct = 32'b11010011100010011100111010111100;
		#400 //-1.7535036e-13 * 1.4813025e-25 = -1183757900000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100111111110111100101001000100;
		b = 32'b11111101001101000011011001000111;
		correct = 32'b10101010001100101101011100010000;
		#400 //2.3780903e+24 * -1.4971429e+37 = -1.588419e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001100100101111010011111110101;
		b = 32'b10110011010101011110010011110110;
		correct = 32'b00011000101101011000001010001100;
		#400 //-2.336632e-31 * -4.9801166e-08 = 4.6919222e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010001101111010111001001010000;
		b = 32'b10101011100001010111001101011101;
		correct = 32'b11100101101101011011010101110100;
		#400 //101708330000.0 * -9.482238e-13 = -1.0726194e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010001011000001111101111010111;
		b = 32'b10110110101010011110000110011001;
		correct = 32'b00011010001010011000010010011000;
		#400 //-1.7748088e-28 * -5.0628555e-06 = 3.505549e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100101010011010001101011010111;
		b = 32'b00101100011110100010101111011010;
		correct = 32'b01111000010100011110001000110000;
		#400 //6.0536265e+22 * 3.555148e-12 = 1.7027776e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010111100111110100010101000101;
		b = 32'b10010011100010101101011001100110;
		correct = 32'b01000011100100101101011010001110;
		#400 //-1.029262e-24 * -3.504751e-27 = 293.6762
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101110010100000101000100101110;
		b = 32'b11001001011000110111111010001101;
		correct = 32'b10100100011010100110101101111001;
		#400 //4.7365827e-11 * -931816.8 = -5.0831695e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110010010100011101011100101101;
		b = 32'b00101000001011110000101011111100;
		correct = 32'b01001001100110010111001000011100;
		#400 //1.2214326e-08 * 9.716833e-15 = 1257027.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010010110110011001101001000011;
		b = 32'b00011101010001111010111110001000;
		correct = 32'b00110101000010110111110000100001;
		#400 //1.3732654e-27 * 2.6428178e-21 = 5.1962166e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101111100101111000000001101100;
		b = 32'b11000101000001001000111011011100;
		correct = 32'b01101010000100100100101011001111;
		#400 //-9.377498e+28 * -2120.9287 = 4.421411e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110001101000111111011011001100;
		b = 32'b11011111000010111001011010111011;
		correct = 32'b01010010000101100101101000000011;
		#400 //-1.6238213e+30 * -1.0058432e+19 = 161438810000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010011000100011011100101011101;
		b = 32'b00111111001011010111111101101110;
		correct = 32'b10010011010101110000010011101110;
		#400 //-1.8392964e-27 * 0.6777257 = -2.7139246e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011000100001001001010001100110;
		b = 32'b11101110010000001000110101111010;
		correct = 32'b00101001101100000100001111111011;
		#400 //-1166183200000000.0 * -1.4898039e+28 = 7.827763e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001001001011011000001011100100;
		b = 32'b10011011110111001001111001100001;
		correct = 32'b10101100110010010101011001111110;
		#400 //2.0885662e-33 * -3.6498297e-22 = -5.722366e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110111100000101011011100101010;
		b = 32'b11111000110101111011000011101100;
		correct = 32'b00111110000110110010010011011000;
		#400 //-5.30245e+33 * -3.4997882e+34 = 0.15150774
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010110101100101110000011000000;
		b = 32'b11010110110001010001110111100100;
		correct = 32'b00111111011010000101000000010101;
		#400 //-98339180000000.0 * -108366085000000.0 = 0.90747195
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110000011101101110100111111;
		b = 32'b00001001100001111011000010011001;
		correct = 32'b01110100000001101100010010010000;
		#400 //0.13951586 * 3.266614e-33 = 4.270963e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001111111000000010110011000110;
		b = 32'b11101110010011000101101011001010;
		correct = 32'b10100001000011000110101000100111;
		#400 //7522061300.0 * -1.5811175e+28 = -4.7574337e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000001100010110011110101110;
		b = 32'b11011010110100011110100000010000;
		correct = 32'b00010100110110000101110010001010;
		#400 //-6.453956e-10 * -2.9541713e+16 = 2.1846927e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010001111101110000011000101110;
		b = 32'b10001011011110111000101110110110;
		correct = 32'b11000101111110110110010111111001;
		#400 //3.8973537e-28 * -4.8445948e-32 = -8044.7466
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010101101000110011111010111000;
		b = 32'b01010110011101101110100010110001;
		correct = 32'b10111110101010010100000101101110;
		#400 //-22436221000000.0 * 67869816000000.0 = -0.3305773
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101101010000101000001110110110;
		b = 32'b11101010011110110101010101111010;
		correct = 32'b00000010010001100010000000110000;
		#400 //-1.1056869e-11 * -7.596101e+25 = 1.455598e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110100000011100101101111101001;
		b = 32'b00101110111000101111000100000101;
		correct = 32'b01000100101000001001011001010110;
		#400 //1.3258217e-07 * 1.0320104e-10 = 1284.698
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111100101010011010001100111000;
		b = 32'b01110100010010100101000000100000;
		correct = 32'b01000111110101101010011101010101;
		#400 //7.046469e+36 * 6.4115545e+31 = 109902.664
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000101100111010000100101111;
		b = 32'b01000100010101000001111110100010;
		correct = 32'b10101011110110001100100011101110;
		#400 //-1.3069775e-09 * 848.49426 = -1.5403492e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011000011100010010010100100001;
		b = 32'b10010110011110111011101011011100;
		correct = 32'b01000001011101010011110001001110;
		#400 //-3.1167265e-24 * -2.0334581e-25 = 15.327223
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110000000111001110110010101;
		b = 32'b01011010001101001101000100000001;
		correct = 32'b00100011001110100101011101100101;
		#400 //0.12853082 * 1.2723825e+16 = 1.0101587e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010110110101010111000011111110;
		b = 32'b10110011110011111111000111100010;
		correct = 32'b01100010100000110110001000100101;
		#400 //-117340640000000.0 * -9.683187e-08 = 1.2117978e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010000111000110000111010111110;
		b = 32'b00101010100111001111010110110001;
		correct = 32'b01100101101110010010101000011101;
		#400 //30475153000.0 * 2.788165e-13 = 1.0930183e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111100101101001110001101111110;
		b = 32'b01110100000100011010010010010101;
		correct = 32'b11001000000111101111100111100100;
		#400 //-7.51382e+36 * 4.6156077e+31 = -162791.56
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001111100110000110100010010111;
		b = 32'b10001011110000101011101011010101;
		correct = 32'b01000011010010000101110011011010;
		#400 //-1.5028644e-29 * -7.5007195e-32 = 200.3627
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010010111001000010110011101110;
		b = 32'b00111110111110110010100001110110;
		correct = 32'b11010011011010001001001100001011;
		#400 //-490003170000.0 * 0.49054307 = -998899400000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111000011111110110010110011001;
		b = 32'b01110011101001100110010110011111;
		correct = 32'b00000100010001000111011001110101;
		#400 //6.0891358e-05 * 2.636665e+31 = 2.3094082e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101100110101111001001011110011;
		b = 32'b11010001100110100010000100100100;
		correct = 32'b11011010101100110000011100100101;
		#400 //2.084904e+27 * -82747620000.0 = -2.5195938e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001001101101011001001011111010;
		b = 32'b11110000111001001111101001001100;
		correct = 32'b00011000010010110000000010001111;
		#400 //-1487455.2 * -5.6692138e+29 = 2.6237417e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011110101001100000000010100111;
		b = 32'b11111110000011101100001011100011;
		correct = 32'b00100000000101001101011010010010;
		#400 //-5.980872e+18 * -4.744057e+37 = 1.2607083e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101000011010101000110011111100;
		b = 32'b00010011001001101100101100011001;
		correct = 32'b11010100101100111111111110000110;
		#400 //-1.30201805e-14 * 2.105228e-27 = -6184689000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100001111100101000010000111011;
		b = 32'b00101110011111111011000110100010;
		correct = 32'b11110010111100101100111010001111;
		#400 //-5.5920503e+20 * 5.8138057e-11 = -9.618571e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111000101011111001101111111011;
		b = 32'b00111001101110000100001010101011;
		correct = 32'b01111110011100111111101100001101;
		#400 //2.8494238e+34 * 0.00035144886 = 8.1076483e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000101000110010100100000000001;
		b = 32'b10110111001101000001001101110011;
		correct = 32'b10001101010110011110100001110110;
		#400 //7.2072505e-36 * -1.0733364e-05 = -6.71481e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011011001010011001000101000101;
		b = 32'b01110011101100011000110100011000;
		correct = 32'b10100110111101000111110100100011;
		#400 //-4.7728997e+16 * 2.8134102e+31 = -1.696482e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000101100011101111011001100001;
		b = 32'b10011100110000100111101000011011;
		correct = 32'b00101000001111000011000001010010;
		#400 //-1.3444121e-35 * -1.2869407e-21 = 1.0446574e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111010100000101000000001100111;
		b = 32'b00001001111001001110010110101001;
		correct = 32'b01110000000100011111010000101100;
		#400 //0.000995648 * 5.5104975e-33 = 1.8068205e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101000010001110111000111100011;
		b = 32'b01011010101101001110101001101011;
		correct = 32'b11001101000011010001110000001111;
		#400 //-3.767407e+24 * 2.546162e+16 = -147964140.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101110010010010011110010001111;
		b = 32'b00101110100110010111110111100111;
		correct = 32'b11111111001001111101000010111010;
		#400 //-1.5569924e+28 * 6.979999e-11 = -2.2306485e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010000110110100000111001101101;
		b = 32'b00001010010001000101011000001010;
		correct = 32'b01000110000011100010100100001111;
		#400 //8.6008065e-29 * 9.453239e-33 = 9098.265
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010111010010101101001001011011;
		b = 32'b01001101110101111110011100011101;
		correct = 32'b10001000111100000111110101010001;
		#400 //-6.5535226e-25 * 452780960.0 = -1.4473936e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100010001001010011110000101100;
		b = 32'b00001101100111000010100010100001;
		correct = 32'b01010100000001110111000010001111;
		#400 //2.2393525e-18 * 9.624023e-31 = 2326836000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000010010011000011010010111100;
		b = 32'b10010101000100100011111100110011;
		correct = 32'b00101100101100101011101001001011;
		#400 //-1.5002687e-37 * -2.953432e-26 = 5.079747e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111101000010110111011100111100;
		b = 32'b10110101001111010101101000001001;
		correct = 32'b11000111001111001000111000011101;
		#400 //0.034049258 * -7.0539005e-07 = -48270.113
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001101001100110001111110101000;
		b = 32'b10011011001000110000000101110000;
		correct = 32'b10110001100011001010100000011100;
		#400 //5.519674e-31 * -1.3483508e-22 = -4.093648e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011010110100000000001100000110;
		b = 32'b01010100000011100111100000000101;
		correct = 32'b10000110001110101110001011110111;
		#400 //-8.603167e-23 * 2447595800000.0 = -3.514946e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100001010010110011011110110101;
		b = 32'b10101001000010111010010110010001;
		correct = 32'b01110111101110100100010011011010;
		#400 //-2.3429395e+20 * -3.1007806e-14 = 7.5559663e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101100001001110010101101010100;
		b = 32'b01100111110011001001010001101100;
		correct = 32'b11000011110100010010111110111111;
		#400 //-8.083809e+26 * 1.9322013e+24 = -418.37302
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011000011001110000111000110110;
		b = 32'b10100001011111010011100100001010;
		correct = 32'b00110110011010011001011011101111;
		#400 //-2.9863225e-24 * -8.5795225e-19 = 3.480756e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111011100110100111100000101000;
		b = 32'b11010111100000010100010111100011;
		correct = 32'b10100011100110001111001011000000;
		#400 //0.004714031 * -284274320000000.0 = -1.6582682e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000110110101001101001111001110;
		b = 32'b01011000010011100100100001111110;
		correct = 32'b10101110000001000000111110001011;
		#400 //-27241.902 * 907243000000000.0 = -3.002713e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111111111001110011111000110111;
		b = 32'b11011110111011111011101110000100;
		correct = 32'b11111111111001110011111000110111;
		#400 //nan * -8.637273e+18 = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100000110001111101000010111010;
		b = 32'b00111110111010011001010101100011;
		correct = 32'b10100001010110101111110110111011;
		#400 //-3.3850035e-19 * 0.45621786 = -7.419708e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100011001001110111111010010111;
		b = 32'b11001100100111101011100100100100;
		correct = 32'b10010110000001110001001011001111;
		#400 //9.0798946e-18 * -83216670.0 = -1.0911148e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001001011110011000110100111110;
		b = 32'b10001010011110001101001011111111;
		correct = 32'b10111110100000000101111111001111;
		#400 //3.0038697e-33 * -1.19804496e-32 = -0.25073096
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111000110000101110110000011001;
		b = 32'b01101011011000011010101111011000;
		correct = 32'b00001100110111010001111001011000;
		#400 //9.2946175e-05 * 2.7281982e+26 = 3.4068704e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111011100100111111100110011110;
		b = 32'b00010011001111110000101110000010;
		correct = 32'b01100111110001100100100101010010;
		#400 //0.0045158407 * 2.4113263e-27 = 1.8727622e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100100011100111011101011111010;
		b = 32'b10011000010101010010100011101011;
		correct = 32'b01001011100100100101101101110101;
		#400 //-5.28506e-17 * -2.7550263e-24 = 19183338.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111111100110110000000010000111;
		b = 32'b10000111010110111100010001111010;
		correct = 32'b01110111101101001000111010001110;
		#400 //-1.2109536 * -1.6533468e-34 = 7.324256e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011100000110111110001101000011;
		b = 32'b10100001111001001111010110000000;
		correct = 32'b00111001101011100100110001111010;
		#400 //-5.1578927e-22 * -1.5514864e-18 = 0.00033244846
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100010110011001010110001101100;
		b = 32'b01011000010010100000011111101111;
		correct = 32'b01001010000000011010110010011010;
		#400 //1.88778e+21 * 888541700000000.0 = 2124582.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101000100101110101000000100110;
		b = 32'b11011010011100101111110100010010;
		correct = 32'b10001101100111110110101001100000;
		#400 //1.6799127e-14 * -1.70988e+16 = -9.82474e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101000010001110100100110010101;
		b = 32'b11101110010000001001000000001000;
		correct = 32'b00111001100001000111100001011001;
		#400 //-3.764433e+24 * -1.4898811e+28 = 0.00025266668
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111001011101010001010011100010;
		b = 32'b11000110101001001110101011000110;
		correct = 32'b00110010001111100011100000110000;
		#400 //-0.000233728 * -21109.387 = 1.1072231e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011111110110011100010100010111;
		b = 32'b10010100101100001110111100101100;
		correct = 32'b01001010100111011000101010110100;
		#400 //-9.222913e-20 * -1.7865795e-26 = 5162330.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101010101110100111111000110000;
		b = 32'b11011010111001101011100000011110;
		correct = 32'b01001111010011101110110101111100;
		#400 //-1.1272805e+26 * -3.2470842e+16 = 3471670300.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101110111010000101100101110101;
		b = 32'b00111011101101011110010111000010;
		correct = 32'b10110010101000111000000010110000;
		#400 //-1.0566029e-10 * 0.005551071 = -1.9034218e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101100101110100001011101011011;
		b = 32'b10110110001110100011111001011011;
		correct = 32'b00110101111111111100101001100101;
		#400 //-5.289031e-12 * -2.7752455e-06 = 1.9057885e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010001111010011000000101001100;
		b = 32'b10001011100000000101100001001100;
		correct = 32'b11000101111010001110000010100111;
		#400 //3.6840604e-28 * -4.943666e-32 = -7452.0815
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010010110110111111000011110001;
		b = 32'b01111011001000100000110110110100;
		correct = 32'b00010111001011011011100100101001;
		#400 //472320080000.0 * 8.4143e+35 = 5.613302e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011010111101100010100110000010;
		b = 32'b10111111110000001111100110000110;
		correct = 32'b10011010101000110100011101111001;
		#400 //1.01810275e-22 * -1.5076149 = -6.753069e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011100011000101100010100100111;
		b = 32'b00011001111000111000011001000111;
		correct = 32'b11000001111111110010011010110100;
		#400 //-7.503194e-22 * 2.3525484e-23 = -31.893898
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001000101100001010111101011010;
		b = 32'b00110101101001001100011001000011;
		correct = 32'b01010010100010010100000010011000;
		#400 //361850.8 * 1.2276654e-06 = 294747100000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100101011101101010110011101110;
		b = 32'b11000101000001010111001101001010;
		correct = 32'b11011111111011001001100111010001;
		#400 //7.280576e+22 * -2135.2056 = -3.4097775e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110101001110110101011000010010;
		b = 32'b01100100100101101010011110101001;
		correct = 32'b10010000000111110010101001010001;
		#400 //-6.978818e-07 * 2.2232742e+22 = -3.138982e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111001100110011000001011111100;
		b = 32'b01111110011011000000100010111011;
		correct = 32'b10111010101001100111111100111111;
		#400 //-9.963476e+34 * 7.8435785e+37 = -0.0012702717
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111101000011111101101111000101;
		b = 32'b00111001001110010010001001100111;
		correct = 32'b11000011010001101110110010101110;
		#400 //-0.035121698 * 0.0001765579 = -198.92453
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111011001001010111101011111100;
		b = 32'b01001000100011010101100000110010;
		correct = 32'b11110010000101011101101101110001;
		#400 //-8.592234e+35 * 289473.56 = -2.9682275e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110100001101110101000011111010;
		b = 32'b01101000010001011000011101111100;
		correct = 32'b00001011011011011001010001110100;
		#400 //1.7072662e-07 * 3.7312218e+24 = 4.5756223e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110101110001110000100100001110;
		b = 32'b01011110010011100001111001000000;
		correct = 32'b11010110111101110011010000000000;
		#400 //-5.046146e+32 * 3.7130947e+18 = -135901355000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010010011001100110110001101001;
		b = 32'b10011010111111011000110000001111;
		correct = 32'b10110110111010001010011100010101;
		#400 //7.270883e-28 * -1.04864624e-22 = -6.9335897e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111000101100101110111001100101;
		b = 32'b01011110000100100010001001001100;
		correct = 32'b10011010000111001011101000110111;
		#400 //-8.532106e-05 * 2.6325156e+18 = -3.2410467e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100000001011110111010010100001;
		b = 32'b01101110000101100010001010101010;
		correct = 32'b10110001100101011001011001001010;
		#400 //-5.057163e+19 * 1.1616164e+28 = -4.3535566e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000101101101111101100110111011;
		b = 32'b11001100101111000011001000001110;
		correct = 32'b10111000011110100001011011101011;
		#400 //5883.2163 * -98668660.0 = -5.962599e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000100011111101111111101000;
		b = 32'b00010100000001000110010100101001;
		correct = 32'b11011100000010110001100100110000;
		#400 //-1.0468257e-09 * 6.684247e-27 = -1.5661086e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011000111110101010101010100000;
		b = 32'b11111000010010110000010000010100;
		correct = 32'b00100000000111100000101100010111;
		#400 //-2204885900000000.0 * -1.6470609e+34 = 1.338679e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100011101001101100100011011010;
		b = 32'b10101000110111001010101100111011;
		correct = 32'b01111010010000010111110100000011;
		#400 //-6.153265e+21 * -2.4499166e-14 = 2.511622e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010111110000010100100111011101;
		b = 32'b00011101111101011001101000001011;
		correct = 32'b10111001010010010111100011010011;
		#400 //-1.2490978e-24 * 6.5010237e-21 = -0.00019213864
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100000101010101010011111110100;
		b = 32'b11111100000000001001100111110101;
		correct = 32'b00100100001010011101101110100110;
		#400 //-9.8376525e+19 * -2.6709465e+36 = 3.6832083e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111100001110011000000000110111;
		b = 32'b00011101010101111111001001001111;
		correct = 32'b11011110010110111110100001000101;
		#400 //-0.011322073 * 2.8580284e-21 = -3.9614978e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010011110000001110000110101011;
		b = 32'b11000010101000011111010000001000;
		correct = 32'b01010000100110000111000110110111;
		#400 //-1656839600000.0 * -80.97662 = 20460714000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111010011010110110100110000100;
		b = 32'b01000001000111010000000011011011;
		correct = 32'b01111000101111111110110010011111;
		#400 //3.0558247e+35 * 9.812709 = 3.1141498e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100010101110011110001111110101;
		b = 32'b01000011010100000100111111001010;
		correct = 32'b01011110111001000111001000101001;
		#400 //1.7145368e+21 * 208.31168 = 8.2306323e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010101100010000000110101111010;
		b = 32'b10000101111010011011001010100000;
		correct = 32'b01001111000101010000100101010011;
		#400 //-5.4951225e-26 * -2.1976831e-35 = 2500416300.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110101000111011001010011010101;
		b = 32'b11101110111011111000111100111101;
		correct = 32'b11000101101010000110010101010111;
		#400 //1.9975812e+32 * -3.707004e+28 = -5388.6675
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000001111111001001111011011110;
		b = 32'b10101110110100101111110010010100;
		correct = 32'b01010010100110010100001000011010;
		#400 //-31.577572 * -9.594561e-11 = 329119500000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011111111010000010101111000011;
		b = 32'b00010110110001010110110100010001;
		correct = 32'b11001000100101101000011011010011;
		#400 //-9.832822e-20 * 3.1895897e-25 = -308278.6
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010110100111000110001101101001;
		b = 32'b01111010000101111001111101111011;
		correct = 32'b00011100000001000000010111011101;
		#400 //85975390000000.0 * 1.9681787e+35 = 4.3682714e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110100101110011110010111001111;
		b = 32'b00111100000010111010100001100111;
		correct = 32'b10111000001010100110000101001010;
		#400 //-3.4626143e-07 * 0.008524037 = -4.0621766e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111110010011110001111100010000;
		b = 32'b11010010111000000010001111011001;
		correct = 32'b11101010111011001000111111101101;
		#400 //6.882787e+37 * -481337050000.0 = -1.4299308e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010100111011001001101100110011;
		b = 32'b10111001100001001000000010010001;
		correct = 32'b00011010111001001001000100010110;
		#400 //-2.3891126e-26 * -0.0002527279 = 9.453299e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111011001111111100101000101011;
		b = 32'b11010011110101100111000100110100;
		correct = 32'b00100110111001001111010100100100;
		#400 //-0.0029264789 * -1842044500000.0 = 1.5887124e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001100100001001101000101000001;
		b = 32'b10000010100111111100111110111111;
		correct = 32'b01001001010101001100001000101100;
		#400 //-2.046376e-31 * -2.348219e-37 = 871458.75
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101101011011101010111111111001;
		b = 32'b11000110010100000001001101100010;
		correct = 32'b11100110100100101101010011000011;
		#400 //4.6168856e+27 * -13316.846 = -3.4669513e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100100101111110101101111001000;
		b = 32'b01010000101111101101001011100010;
		correct = 32'b11010011100000000101101111010100;
		#400 //-2.8239533e+22 * 25611932000.0 = -1102592900000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101111111010110100100101100010;
		b = 32'b01110000010110001001100011101100;
		correct = 32'b00111111000010110000101101101011;
		#400 //1.4563538e+29 * 2.6813453e+29 = 0.543143
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111101101000111010101110001100;
		b = 32'b00010111010001001001101111111000;
		correct = 32'b11100101110101010001110001011011;
		#400 //-0.07991704 * 6.3527876e-25 = -1.2579839e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101110011001100000001011011111;
		b = 32'b01001001110011111101000101100001;
		correct = 32'b11100100000011011010101101011110;
		#400 //-1.7796256e+28 * 1702444.1 = -1.0453357e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011010101000010000011011011110;
		b = 32'b11010100100011001011011101010001;
		correct = 32'b01000101100100100111100110101111;
		#400 //-2.266251e+16 * -4834967700000.0 = 4687.2104
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010110100011000101000100001010;
		b = 32'b11011001010010000100001011111110;
		correct = 32'b00111100101100110101111011011001;
		#400 //-77139840000000.0 * -3523041000000000.0 = 0.021895813
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111011100011001010011011101010;
		b = 32'b11111110001100110011111000000000;
		correct = 32'b10111100110010001110001001011000;
		#400 //1.460614e+36 * -5.9563433e+37 = -0.024521992
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001101000001011101000111001100;
		b = 32'b11000010101111111000101100111000;
		correct = 32'b11001001101100101101100111011001;
		#400 //140319940.0 * -95.77191 = -1465147.1
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101000110111110010100111011111;
		b = 32'b10110111100000010110111010100011;
		correct = 32'b11110000110111001011000110111010;
		#400 //8.430881e+24 * -1.5429518e-05 = -5.464125e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010001010110111001011100100110;
		b = 32'b11010110000011001011110110110010;
		correct = 32'b10111010110001111011011000011011;
		#400 //58945855000.0 * -38686590000000.0 = -0.0015236767
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110001010001010110001011011011;
		b = 32'b01100000000001010110011110000101;
		correct = 32'b01010000101111010110001111001010;
		#400 //9.774089e+29 * 3.8451193e+19 = 25419469000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000100011011011001100001111000;
		b = 32'b10100111001110011000111111111110;
		correct = 32'b10011100101000111110010001100101;
		#400 //2.7929226e-36 * -2.5751966e-15 = -1.0845474e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110000111101001000001111010;
		b = 32'b01010111010100011100111011111101;
		correct = 32'b10011110010000010111100101010001;
		#400 //-2.362793e-06 * 230686940000000.0 = -1.02424226e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001100001010111001000011100100;
		b = 32'b00001100100000110010010011011011;
		correct = 32'b01111111001001110111001111110101;
		#400 //44974990.0 * 2.0205927e-31 = 2.2258316e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010110010111001100001100001111;
		b = 32'b11000110011100111111111011111000;
		correct = 32'b10001111011001111001111101110111;
		#400 //1.7833008e-25 * -15615.742 = -1.1419891e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001110001100010101001001001011;
		b = 32'b01110100011011111101000010110000;
		correct = 32'b00011001001111010100100111100101;
		#400 //743740100.0 * 7.6000466e+31 = 9.785994e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010100000100011001011111010001;
		b = 32'b10111100100010001110010001010001;
		correct = 32'b10010111000010000010001011010000;
		#400 //7.35057e-27 * -0.016710432 = -4.398791e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110101000101100000000110110101;
		b = 32'b11101101110100101001001001000111;
		correct = 32'b10000110101101100101111001111011;
		#400 //5.588184e-07 * -8.1460863e+27 = -6.859962e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111100010111111000111001011010;
		b = 32'b10001000111001110000110101000100;
		correct = 32'b11110010111101111011000111100011;
		#400 //0.013644779 * -1.39059255e-33 = -9.812205e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001010100111001100001100011101;
		b = 32'b00011110011101010101111000110001;
		correct = 32'b11101011101000111000111000001010;
		#400 //-5136782.5 * 1.298967e-20 = -3.9545134e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010100010000111110010001001101;
		b = 32'b00111100001100110101000001001010;
		correct = 32'b11010111100010111101010110000100;
		#400 //-3365395500000.0 * 0.010944435 = -307498320000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011111110001010001011100101100;
		b = 32'b01000110100111000010001010010010;
		correct = 32'b11011000101000011001001101001111;
		#400 //-2.8403737e+19 * 19985.285 = -1421232500000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011100010000101100110111001110;
		b = 32'b01110011111101101101010101101010;
		correct = 32'b10100111110010100000100111000010;
		#400 //-2.1932972e+17 * 3.9112353e+31 = -5.6076842e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111100101001111000001001000100;
		b = 32'b01101000101010101000011010111111;
		correct = 32'b01010011011110110111100001010011;
		#400 //6.9580454e+36 * 6.4423034e+24 = 1080055500000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101011011111001010001101111011;
		b = 32'b10011111011011001011001000000010;
		correct = 32'b11001011100010001001111100101101;
		#400 //8.975526e-13 * -5.012219e-20 = -17907290.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110000101110010011101011110000;
		b = 32'b11111111110001111101100100011100;
		correct = 32'b11111111110001111101100100011100;
		#400 //-4.5860782e+29 * nan = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110101010111001110101011111011;
		b = 32'b11011011111101011110101011011011;
		correct = 32'b01011000111001011111100110111011;
		#400 //-2.800467e+32 * -1.3843919e+17 = 2022886000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111000011110000000001001110101;
		b = 32'b10111110001110010110111001110111;
		correct = 32'b00111001101010110011001001001111;
		#400 //-5.9130096e-05 * -0.18108545 = 0.00032653144
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101011011111010000100000100000;
		b = 32'b10111100000111101000000000011001;
		correct = 32'b00101110110011000101011100110001;
		#400 //-8.989493e-13 * -0.009674096 = 9.292334e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000000011111111010100100011101;
		b = 32'b00101110110100101100110100001011;
		correct = 32'b01010001000110110011110100111000;
		#400 //3.9946969 * 9.586117e-11 = 41671690000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001001110011000001000000001101;
		b = 32'b01010110011011000000111110001011;
		correct = 32'b10110010110111010100110010011001;
		#400 //-1671681.6 * 64887875000000.0 = -2.5762619e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011110001000010011100111011011;
		b = 32'b01111001000110100100000111001111;
		correct = 32'b10100100100001011100100001011111;
		#400 //-2.9043894e+18 * 5.005928e+34 = -5.8019e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001101010101110000000101000100;
		b = 32'b11101010111101011001100001000101;
		correct = 32'b10100001111000000001110100111000;
		#400 //225449020.0 * -1.4845295e+26 = -1.5186565e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101101000000011110001000000111;
		b = 32'b11001111110000001110000000110010;
		correct = 32'b11011100101011000110010000010010;
		#400 //2.512301e+27 * -6471836700.0 = -3.881898e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010111000110100100100101000100;
		b = 32'b01111111111010110000001001010111;
		correct = 32'b01111111111010110000001001010111;
		#400 //169639460000000.0 * nan = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011000001101110101011100001100;
		b = 32'b10100101000110010100010000001001;
		correct = 32'b11110010100110010001110111010110;
		#400 //806337970000000.0 * -1.3293686e-16 = -6.0655713e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000110110001100111010100101100;
		b = 32'b01110100011010010011010101111011;
		correct = 32'b10010001110110011101101001000101;
		#400 //-25402.586 * 7.3906853e+31 = -3.4371082e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110100100101101110000100010000;
		b = 32'b10101100111000101100111011011101;
		correct = 32'b01000111001010100100110001101000;
		#400 //-2.8103432e-07 * -6.4462728e-12 = 43596.406
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010110100110011100010111011000;
		b = 32'b10100100111101100100001100000111;
		correct = 32'b01110001000111111101101010000111;
		#400 //-84537506000000.0 * -1.0679904e-16 = 7.915568e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000001111100110001111100000010;
		b = 32'b00011100000000110010100100101100;
		correct = 32'b10100101011011010100001100011110;
		#400 //-8.9308596e-38 * 4.339748e-22 = -2.0579213e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001011011000100111110000110101;
		b = 32'b11000101001001011011000111101010;
		correct = 32'b11000101101011101111010111101110;
		#400 //14842933.0 * -2651.1196 = -5598.741
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101010001011111100011001110010;
		b = 32'b00111010010001010101000111110010;
		correct = 32'b11101111011001000000110001000111;
		#400 //-5.3124787e+25 * 0.00075271644 = -7.0577425e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101001001101100011010001000011;
		b = 32'b11011101010000111110110000000011;
		correct = 32'b01001011011011100001001101100110;
		#400 //-1.3766956e+25 * -8.823539e+17 = 15602534.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111001010110110000001011000011;
		b = 32'b11111100101011001100011000001110;
		correct = 32'b00111100001000100100000101000101;
		#400 //-7.1073064e+34 * -7.176737e+36 = 0.009903257
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111100001011000000001001101;
		b = 32'b11111111001111110000100001000110;
		correct = 32'b10000111101100101110011100111011;
		#400 //68352.6 * -2.539255e+38 = -2.6918368e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111010100101110101110011110101;
		b = 32'b00100101100001001000101100001001;
		correct = 32'b01010100100100100010110011001000;
		#400 //0.0011548089 * 2.2992564e-16 = 5022532000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011101001010010111001110110011;
		b = 32'b10011110100110111011101101010111;
		correct = 32'b00111110000010110100011011100110;
		#400 //-2.2426779e-21 * -1.6488745e-20 = 0.13601264
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111001011100101001100011110000;
		b = 32'b11101100001000100110011110011001;
		correct = 32'b00001100101111110011010001001011;
		#400 //-0.00023135892 * -7.853408e+26 = 2.9459682e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000010011110100100011110110100;
		b = 32'b01111110010010100000110001111000;
		correct = 32'b00000011100111101000111000011011;
		#400 //62.570023 * 6.71422e+37 = 9.319031e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000000011000100101100010100101;
		b = 32'b10011011011011110110101001110100;
		correct = 32'b10100100010100100101000100111010;
		#400 //9.031678e-39 * -1.9804013e-22 = -4.5605293e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110010110001010010001010010111;
		b = 32'b01101101011001000101110000000011;
		correct = 32'b11000100110111001111111100001110;
		#400 //-7.8093265e+30 * 4.4171136e+27 = -1767.9705
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100100010011101100001011010101;
		b = 32'b11110111100001010011010101011101;
		correct = 32'b00101100010001101010110100111101;
		#400 //-1.5256274e+22 * -5.403577e+33 = 2.8233659e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110100011010010100000001010100;
		b = 32'b11110001101000001000101101111000;
		correct = 32'b11000010001110011111011111000010;
		#400 //7.392028e+31 * -1.5899587e+30 = -46.49195
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111100100110010101011001100100;
		b = 32'b01111001110110100111000110011001;
		correct = 32'b11000010001100111011001101000010;
		#400 //-6.369389e+36 * 1.4177809e+35 = -44.925056
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101010111100010101011110111010;
		b = 32'b00111000111100110011111011100110;
		correct = 32'b10110001011111011111111101001001;
		#400 //-4.2871072e-13 * 0.00011598859 = -3.6961458e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001111010101101100110101110000;
		b = 32'b00111111100000001101101001000110;
		correct = 32'b11001111010101010110000110010001;
		#400 //-3603787800.0 * 1.0066612 = -3579941000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100010010000111111101000110011;
		b = 32'b10000011111011101001100011100111;
		correct = 32'b01011101110100100100010101111111;
		#400 //-2.6559882e-18 * -1.4023487e-36 = 1.893957e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001111111110010001110111101110;
		b = 32'b00110001100011111011001011000111;
		correct = 32'b01011101110111011110011011110000;
		#400 //8358976500.0 * 4.1821724e-09 = 1.9987164e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110111001100000111111101010000;
		b = 32'b01111101100011110000110110110101;
		correct = 32'b10111001000111011110110010101011;
		#400 //-3.5797908e+33 * 2.3768847e+37 = -0.00015060852
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111100101100011011000111111111;
		b = 32'b00111101000010000010010011001010;
		correct = 32'b00111111001001110001000011101100;
		#400 //0.02169132 * 0.03323821 = 0.65260196
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111011110110000110010010000011;
		b = 32'b01111000001010010110010111101001;
		correct = 32'b00000011001000111000001010000110;
		#400 //0.006603779 * 1.3743206e+34 = 4.805123e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110101100001101001101001001111;
		b = 32'b01110010001111101100010110101001;
		correct = 32'b11000010101101001010000000100001;
		#400 //-3.4125856e+32 * 3.778631e+30 = -90.31275
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000001010011111100100010100010;
		b = 32'b01100111110011111100010010011100;
		correct = 32'b10011001000000000000001001111011;
		#400 //-12.986483 * 1.9623133e+24 = -6.617946e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011111110111011001111011100011;
		b = 32'b10010000000000011001101000100101;
		correct = 32'b11001111010110101110000110001001;
		#400 //9.3859997e-20 * -2.5559513e-29 = -3672213800.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001000010010000011001001110010;
		b = 32'b10010111011111100101101100010111;
		correct = 32'b10110000010010010111110110111100;
		#400 //6.024461e-34 * -8.21868e-25 = -7.3302053e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011010011111001101110100001000;
		b = 32'b11001100011100001001010001101010;
		correct = 32'b01001101100001101000100100010110;
		#400 //-1.779368e+16 * -63066536.0 = 282141380.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010010110010101000011000101000;
		b = 32'b00101001110011111111011011001001;
		correct = 32'b01101000011110010100110110110011;
		#400 //434917080000.0 * 9.235457e-14 = 4.7092102e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001010011001000001001110000011;
		b = 32'b01011001100110101000111101001001;
		correct = 32'b10110000001111001110001000100011;
		#400 //-3736800.8 * 5438086000000000.0 = -6.871536e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010010101101100100100000001111;
		b = 32'b11110000111011010110010101100101;
		correct = 32'b10100001010001001001000011110111;
		#400 //391446500000.0 * -5.877642e+29 = -6.659924e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001000111111111101011111010110;
		b = 32'b11111011000010000000101010001101;
		correct = 32'b10001101011100001011100001110111;
		#400 //523966.7 * -7.063664e+35 = -7.417775e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011101000001001010011011110100;
		b = 32'b11001011000011110110100001010001;
		correct = 32'b01010001011011001100110011101000;
		#400 //-5.974122e+17 * -9398353.0 = 63565627000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101000110001111101110001100111;
		b = 32'b00001001101000000010001110110101;
		correct = 32'b01011110100111111011111111011111;
		#400 //2.2189022e-14 * 3.8552178e-33 = 5.755582e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101000000001010101100101111010;
		b = 32'b00111000010010111110100110111100;
		correct = 32'b00101111001001110110100101110101;
		#400 //7.402385e-15 * 4.8616654e-05 = 1.5226027e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101011111111001000111001011000;
		b = 32'b00011110010010100100110010001011;
		correct = 32'b01001101000111111100110010001010;
		#400 //1.7945185e-12 * 1.070962e-20 = 167561380.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101011010100010111111110110000;
		b = 32'b00110101111011010000001010011111;
		correct = 32'b00110100111000100100100011000110;
		#400 //7.442892e-13 * 1.7658639e-06 = 4.214873e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100011010001001100110001100001;
		b = 32'b11110011101110001101000010011110;
		correct = 32'b00101111000010000100110010101111;
		#400 //-3.630289e+21 * -2.9285092e+31 = 1.2396371e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101100111011101000111001001101;
		b = 32'b00111010010010000011011111011011;
		correct = 32'b01110010000110001000001001100110;
		#400 //2.3071707e+27 * 0.00076377176 = 3.0207593e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001101111110100001110000110000;
		b = 32'b01110111110110001000101101101111;
		correct = 32'b10010101100100111101011100110010;
		#400 //-524518900.0 * 8.784095e+33 = -5.9712346e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000101011111111110101110110001;
		b = 32'b10000110000011101100101111100101;
		correct = 32'b10111110111001010110011100000001;
		#400 //1.2033332e-35 * -2.685703e-35 = -0.44805148
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001010011100111111010100101011;
		b = 32'b01101100011110011001100111110001;
		correct = 32'b00011101011110100011011000110000;
		#400 //3997002.8 * 1.206998e+27 = 3.3115239e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000101111000011100010110011100;
		b = 32'b00110001101111100110110111000101;
		correct = 32'b00010011100101111100000110101001;
		#400 //2.1231489e-35 * 5.542207e-09 = 3.8308723e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010000101100100110110001111101;
		b = 32'b00101001010001111010111100100000;
		correct = 32'b00100110111001001011111001100111;
		#400 //7.0375773e-29 * 4.4338773e-14 = 1.5872287e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111111110001110101010001111110;
		b = 32'b11101010100011011111100100000111;
		correct = 32'b00010100101100111011011001010111;
		#400 //-1.557266 * -8.581727e+25 = 1.8146301e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010110100011100011011100000111;
		b = 32'b10101011011000001101100100000011;
		correct = 32'b00101010101000011110101100101010;
		#400 //-2.2976064e-25 * -7.988195e-13 = 2.8762523e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110111111110100101111010111001;
		b = 32'b01100111110011100110000010000101;
		correct = 32'b11001111100110110100100100010111;
		#400 //-1.0156214e+34 * 1.949176e+24 = -5210517000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011011100110110001110000001101;
		b = 32'b01111000111001101100000110111111;
		correct = 32'b10100010001011000001001111010101;
		#400 //-8.731893e+16 * 3.7442435e+34 = -2.3320846e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000100101101011111101100011111;
		b = 32'b11001101001001111101111001101011;
		correct = 32'b00110111000010101100001010110000;
		#400 //-1455.8475 * -176023220.0 = 8.27077e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101100110100001111100011010000;
		b = 32'b00111010000010111001010111011110;
		correct = 32'b01110010001111111010000010100101;
		#400 //2.0210524e+27 * 0.0005324761 = 3.795574e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111101000010011100110001111101;
		b = 32'b10001000001110110101111101110000;
		correct = 32'b01110100001111000100010011011101;
		#400 //-0.03364228 * -5.638545e-34 = 5.9664827e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010001010100011001000010101111;
		b = 32'b11100101010101000110011011011010;
		correct = 32'b10101011011111001001010011000111;
		#400 //56254722000.0 * -6.2689936e+22 = -8.9734855e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110011100110010000111011000100;
		b = 32'b10000001010111101000111100011010;
		correct = 32'b11110001101100000000111000111110;
		#400 //7.1273035e-08 * -4.087763e-38 = -1.7435705e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000110110100010111100001110100;
		b = 32'b10000000110100110010111011110111;
		correct = 32'b11000101011111011110110001101110;
		#400 //7.879405e-35 * -1.9394138e-38 = -4062.7769
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011101010100110111001011000001;
		b = 32'b00101011110010001101111110001100;
		correct = 32'b10110001000001101011110100010101;
		#400 //-2.7984944e-21 * 1.4272901e-12 = -1.9607047e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100101011011111011000010011101;
		b = 32'b01100010010110100111100001001100;
		correct = 32'b11000010100011000110111011000010;
		#400 //-7.074397e+22 * 1.0075146e+21 = -70.216324
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110100111101011100110110001011;
		b = 32'b11101010111000110001011111101101;
		correct = 32'b11001001100010101000101110100100;
		#400 //1.557961e+32 * -1.3726957e+26 = -1134964.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110001001111110001011111101001;
		b = 32'b10111100100011011110110001011110;
		correct = 32'b00110100001011000101100010100110;
		#400 //-2.780775e-09 * -0.017324623 = 1.6050998e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100101111010100100101000010;
		b = 32'b10011010010100110101001011010000;
		correct = 32'b11101001111001010100110110111111;
		#400 //1514.2893 * -4.3700673e-23 = -3.4651395e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101011101111111111101001010110;
		b = 32'b11100000101010010101001110111001;
		correct = 32'b00001010100100010001111101011110;
		#400 //-1.3640848e-12 * -9.761039e+19 = 1.3974791e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010100011001111111101000110111;
		b = 32'b11001010011011011111001100010001;
		correct = 32'b11001001011110011001001100101100;
		#400 //3985341400000.0 * -3898564.2 = -1022258.75
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101011001100100000000100111111;
		b = 32'b11100000100101110010001001000011;
		correct = 32'b00001010000101101100001000000111;
		#400 //-6.3240033e-13 * -8.712272e+19 = 7.25873e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010010001101100011100100000011;
		b = 32'b00000111010110111101110000010111;
		correct = 32'b01001010010101000010110100011111;
		#400 //5.7499346e-28 * 1.6540407e-34 = 3476295.8
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111101111111000100110010101100;
		b = 32'b01110001001110110001101010101010;
		correct = 32'b10001100001011001001100111010001;
		#400 //-0.123193115 * 9.264949e+29 = -1.3296685e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010100110010011000110110001100;
		b = 32'b00000100110110101111011100110111;
		correct = 32'b01001111011010111010010001100101;
		#400 //2.0351644e-26 * 5.1478585e-36 = 3953419500.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000101101110101011101011111011;
		b = 32'b10001100001111110101110100100010;
		correct = 32'b11111000111110011100110100110101;
		#400 //5975.3726 * -1.4742131e-31 = -4.0532625e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100110100111010101000001100011;
		b = 32'b10111000101100100010111011100011;
		correct = 32'b10101101011000100000010001001101;
		#400 //1.0915852e-15 * -8.496435e-05 = -1.2847568e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011011001100011111110000111000;
		b = 32'b01001001011100000100111100101011;
		correct = 32'b01010001001111011001101101001010;
		#400 //5.009839e+16 * 984306.7 = 50897134000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110000100110110000001010011010;
		b = 32'b01011101011000010000111011001110;
		correct = 32'b00010010101100000101001001100001;
		#400 //1.1278474e-09 * 1.01357036e+18 = 1.11274695e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010010010101100011001111000110;
		b = 32'b10011000011011101111111110110010;
		correct = 32'b10111001011001010111000010000101;
		#400 //6.759031e-28 * -3.0889872e-24 = -0.00021881059
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111010110110100101010100011100;
		b = 32'b11111000111010010010101111100110;
		correct = 32'b10000001011011111011010101001011;
		#400 //0.0016657445 * -3.7834235e+34 = -4.4027438e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100100110111011001111101010101;
		b = 32'b01101000100111000101100011111110;
		correct = 32'b00111011101101010111000010010000;
		#400 //3.2705692e+22 * 5.9066463e+24 = 0.0055371
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011100010000101101010110001;
		b = 32'b11001110100110011111111010001100;
		correct = 32'b00111100011000101010110011011001;
		#400 //-17872226.0 * -1291798000.0 = 0.013835155
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110101011110010110100000111000;
		b = 32'b01101011101001010010111000110110;
		correct = 32'b01001001010000010100010010011101;
		#400 //3.1616107e+32 * 3.9938197e+26 = 791625.8
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011100001100011100111110010000;
		b = 32'b01000001000010110001011111010110;
		correct = 32'b10011010101000111010000100111100;
		#400 //-5.8832656e-22 * 8.693319 = -6.767571e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010110110011101110000110001010;
		b = 32'b00110110010001100001101100101000;
		correct = 32'b10100000000001011010101101101110;
		#400 //-3.342343e-25 * 2.9520106e-06 = -1.132226e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000001111101111010110101111001;
		b = 32'b00111001101000010100110000000100;
		correct = 32'b11000111110001001000110010000101;
		#400 //-30.959703 * 0.0003076495 = -100633.04
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001101010111010100111111110110;
		b = 32'b10011110111001000110000101111011;
		correct = 32'b00101101111110000001001110100101;
		#400 //-6.819713e-31 * -2.4180756e-20 = 2.820306e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011000111111111000100110001110;
		b = 32'b10001011111110100001001111101110;
		correct = 32'b01001100100000101100101101011100;
		#400 //-6.605485e-24 * -9.6326484e-32 = 68573920.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010110101110010000011011011101;
		b = 32'b11000100010111111110110110110000;
		correct = 32'b10010001110100111000011011011010;
		#400 //2.9892693e-25 * -895.71387 = -3.337304e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000110110110110000110111100000;
		b = 32'b11010100001000011001110001100010;
		correct = 32'b00110010001011010111111100100010;
		#400 //-28038.938 * -2776453600000.0 = 1.0098832e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101001000100101000111111111000;
		b = 32'b00111001101101101000000101001010;
		correct = 32'b10101110110011011001010101001100;
		#400 //-3.2543385e-14 * 0.00034810073 = -9.348841e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110100001001011000001001111000;
		b = 32'b00011011111100101010011110111001;
		correct = 32'b01010111101011101001110010100011;
		#400 //1.5414287e-07 * 4.014393e-22 = 383975550000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101110000101011011111101101000;
		b = 32'b10010010111111101111011111000000;
		correct = 32'b11011010100101100101101010011011;
		#400 //3.404868e-11 * -1.6090729e-27 = -2.1160434e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010011000010110000101110101010;
		b = 32'b11110111001010110011110011110110;
		correct = 32'b00011011010011111101111101001111;
		#400 //-597196140000.0 * -3.473122e+33 = 1.7194794e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000001011111110000100101011110;
		b = 32'b01101101110010011000100100000001;
		correct = 32'b00010011001000011111101011100111;
		#400 //15.939787 * 7.7965143e+27 = 2.0444761e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011000100001111100100101101011;
		b = 32'b10110110101001110110010011000001;
		correct = 32'b10100001010011111010100110101101;
		#400 //3.5100062e-24 * -4.988717e-06 = -7.035889e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001101101011010110011111000010;
		b = 32'b01110001110110011100111100101001;
		correct = 32'b00011011010010111100111101101110;
		#400 //363657280.0 * 2.157078e+30 = 1.685879e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000101101010010100001011001000;
		b = 32'b01001101111111110110011110010111;
		correct = 32'b10110111001010011010011111001001;
		#400 //-5416.3477 * 535622370.0 = -1.01122505e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101110111001101111010001001011;
		b = 32'b01010010000100010001101110010010;
		correct = 32'b01011100010010111011100110111110;
		#400 //3.5738442e+28 * 155808200000.0 = 2.2937458e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100000111001010111011100000101;
		b = 32'b11011100001110000010000001100001;
		correct = 32'b00000100000111111000010010100011;
		#400 //-3.887287e-19 * -2.0730799e+17 = 1.8751264e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001110110011110111001100110011;
		b = 32'b11101000001101100101101011010101;
		correct = 32'b10100110000100011001110101110010;
		#400 //1740216700.0 * -3.444585e+24 = -5.052036e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000100111100001111111011011;
		b = 32'b10010110000100100101010011101010;
		correct = 32'b01011010000010100101000010111110;
		#400 //-1.1505067e-09 * -1.182058e-25 = 9733081000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101011101110110010110000000101;
		b = 32'b11001000100010110000100010010001;
		correct = 32'b01100010101011000101000101111100;
		#400 //-4.52554e+26 * -284740.53 = 1.5893558e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000110001110111000010111110100;
		b = 32'b10111010001101100000000111101000;
		correct = 32'b11001011100000111110000100001100;
		#400 //12001.488 * -0.0006943033 = -17285656.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101001001000000001001101100100;
		b = 32'b01100001100100010000000100000101;
		correct = 32'b01000111000011010100110111101011;
		#400 //1.2094981e+25 * 3.3435642e+20 = 36173.918
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001110111111100101111101001111;
		b = 32'b00111001101010111000110111010100;
		correct = 32'b00010100101111011100101011011101;
		#400 //6.2707613e-30 * 0.00032721332 = 1.9164138e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000001010011001001000010010011;
		b = 32'b10101011010101001101001111110100;
		correct = 32'b01010101011101100000111110000100;
		#400 //-12.785296 * -7.5611674e-13 = 16909156000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010100100101011110010000110001;
		b = 32'b11001010101100101100010101110010;
		correct = 32'b01001001010101101010010011100001;
		#400 //-5150228300000.0 * -5857977.0 = 879182.06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110101010110101101111101011111;
		b = 32'b01100000001001010011000111110101;
		correct = 32'b11010100101010011001011101101010;
		#400 //-2.7745391e+32 * 4.761426e+19 = -5827118000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110010011100100111011110111011;
		b = 32'b11000010101101110010010100101110;
		correct = 32'b11101111001010010111010111011101;
		#400 //4.8025675e+30 * -91.57262 = -5.2445455e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001111011101000010010110000111;
		b = 32'b11101010011111000010010001000000;
		correct = 32'b00100100011101111110000111110101;
		#400 //-4096100000.0 * -7.6205123e+25 = 5.375098e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010111100010110100111100000100;
		b = 32'b01101101111010000011100110111001;
		correct = 32'b10101001000110011001001000010110;
		#400 //-306342970000000.0 * 8.983788e+27 = -3.4099534e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101000010111001000101111011111;
		b = 32'b11011100111110100111110000110001;
		correct = 32'b10001010111000010110011011110000;
		#400 //1.2242783e-14 * -5.6404235e+17 = -2.1705433e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001001111100001010010000101111;
		b = 32'b11010100100100000111001001001010;
		correct = 32'b10110100110101010011111000001000;
		#400 //1971333.9 * -4963142000000.0 = -3.9719475e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100111010100110010101101010000;
		b = 32'b10111111100100110001101110110000;
		correct = 32'b10100111001101111011110101110010;
		#400 //2.9305612e-15 * -1.1492825 = -2.549905e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110111100001011000000110001100;
		b = 32'b01001100100101101110110101111110;
		correct = 32'b00101010011000100111001100100101;
		#400 //1.591516e-05 * 79129580.0 = 2.0112781e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110110011001011111011100011110;
		b = 32'b11010010001001011110011100000010;
		correct = 32'b01100011101100010110110101001111;
		#400 //-1.1660626e+33 * -178136320000.0 = 6.5459004e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010101010011110010011110110000;
		b = 32'b10000000010010111000111110010101;
		correct = 32'b11010100101011110111010111001101;
		#400 //4.1834625e-26 * -6.93917e-39 = -6028765000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111001000001011111111110111111;
		b = 32'b00000011110010110111001101110000;
		correct = 32'b01110100101010001001110000000100;
		#400 //0.00012779141 * 1.1957771e-36 = 1.0686893e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111111111111000010011101101100;
		b = 32'b11101000111101111110010110100001;
		correct = 32'b01111111111111000010011101101100;
		#400 //nan * -9.3652834e+24 = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001001001111101111010100011000;
		b = 32'b10101000110110110101100111011111;
		correct = 32'b10011111110111101101110011000011;
		#400 //2.298566e-33 * -2.435286e-14 = -9.438588e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001000001101111111000010010000;
		b = 32'b01101111001101110010010110000000;
		correct = 32'b10011000100000001000110111101011;
		#400 //-188354.25 * 5.668109e+28 = -3.3230525e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101010001010011001011111111011;
		b = 32'b01010110110110101110000111000010;
		correct = 32'b11010010110001100101101001111110;
		#400 //-5.1256543e+25 * 120331580000000.0 = -425960870000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110011101110000011010000011100;
		b = 32'b01000011111001010010111101011001;
		correct = 32'b11101111010011011100000101110101;
		#400 //-2.9188218e+31 * 458.3699 = -6.36783e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001010100011010010011001110010;
		b = 32'b11100011110101110111010100100011;
		correct = 32'b00100110001001111011010111010100;
		#400 //-4625209.0 * -7.948981e+21 = 5.8186187e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101110001101011000011001100000;
		b = 32'b10000000001001001010111111001000;
		correct = 32'b01101110000111100101010111100001;
		#400 //-4.1273984e-11 * -3.369136e-39 = 1.2250613e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101000001101111011101011000111;
		b = 32'b11101110001010011000010010110111;
		correct = 32'b10111001100010101011101100000111;
		#400 //3.470554e+24 * -1.3115852e+28 = -0.00026460757
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100000011011000101000011110001;
		b = 32'b11011001100101100011000011110110;
		correct = 32'b01000110010010010110011001010010;
		#400 //-6.81135e+19 * -5284385000000000.0 = 12889.58
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011100010011001101000110111101;
		b = 32'b11000111101000110001010011000000;
		correct = 32'b11010100001000001100001001111111;
		#400 //2.3060602e+17 * -83497.5 = -2761831500000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000110100110010111100000101000;
		b = 32'b00100101110011101100000100111110;
		correct = 32'b00100000001111100000010111011101;
		#400 //5.772876e-35 * 3.586625e-16 = 1.6095566e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100001110000101101001011111001;
		b = 32'b11100111011101010000001100101001;
		correct = 32'b00111001110010111000111110100010;
		#400 //-4.492338e+20 * -1.1570381e+24 = 0.00038826192
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110001011011011111111001100010;
		b = 32'b11110100010011100110111101100010;
		correct = 32'b00111100100100111001000101100010;
		#400 //-1.1784876e+30 * -6.542189e+31 = 0.01801366
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001101110110000100000010101010;
		b = 32'b11010010000111111001110111001011;
		correct = 32'b10111011001011010110101011111001;
		#400 //453514560.0 * -171386780000.0 = -0.0026461466
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000100101100100101000010110010;
		b = 32'b10100010110101101000011000000010;
		correct = 32'b10100001010101001100101010001001;
		#400 //4.1921706e-36 * -5.8146703e-18 = -7.2096447e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000100100100100011111010101101;
		b = 32'b00000100101100010001101000100010;
		correct = 32'b10111111010100110110010101100010;
		#400 //-3.4381994e-36 * 4.16365e-36 = -0.8257657
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001100111101010011010010010100;
		b = 32'b00101111000011011000101011010011;
		correct = 32'b10011101010111011011111010110110;
		#400 //-3.7779871e-31 * 1.2873196e-10 = -2.9347702e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011110101000000100100111101001;
		b = 32'b10010101100100111010010101111001;
		correct = 32'b11001000100010101111010111001001;
		#400 //1.6971227e-20 * -5.96339e-26 = -284590.28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100001000100111111000111001010;
		b = 32'b01010011111011100100100111100110;
		correct = 32'b00001100100111101111000011011000;
		#400 //5.012554e-19 * 2046884000000.0 = 2.4488707e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011000011011101011000111100011;
		b = 32'b10111110101101011000100011101000;
		correct = 32'b11011001001010000100110110110011;
		#400 //1049791140000000.0 * -0.35456014 = -2960826700000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011000110001101011010111110000;
		b = 32'b11101101011101011000011001101111;
		correct = 32'b00101010110011110011000000110101;
		#400 //-1747877700000000.0 * -4.7491467e+27 = 3.6804037e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011001111000010010000001011001;
		b = 32'b11001000111110000110001010110000;
		correct = 32'b11010000011010000000011100100000;
		#400 //7920929500000000.0 * -508693.5 = -15571124000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110101110010101111100010110;
		b = 32'b01010000001011111100111100011111;
		correct = 32'b00101110000001101111011001000110;
		#400 //0.36205357 * 11798347000.0 = 3.0686807e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000100110000100000111100010000;
		b = 32'b00100100010000001010110100101100;
		correct = 32'b00100000000000001110101100011001;
		#400 //4.5623014e-36 * 4.1780046e-17 = 1.0919809e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010010101100111010100101011110;
		b = 32'b10011001110101101010000110010110;
		correct = 32'b10111000010101100100101001001100;
		#400 //1.133824e-27 * -2.2192345e-23 = -5.109077e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001100000011111010000110110001;
		b = 32'b10010111001100011110000111101010;
		correct = 32'b00110100010011101011010100110001;
		#400 //-1.1064977e-31 * -5.747693e-25 = 1.9251162e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100000001010101101000011110001;
		b = 32'b01111011000110100001100100000111;
		correct = 32'b10100100100011011110001100010011;
		#400 //-4.923441e+19 * 8.001213e+35 = -6.153368e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111000100001100001011100111100;
		b = 32'b10000010001011101000011110100111;
		correct = 32'b11110101110001001010111100011010;
		#400 //6.393946e-05 * -1.2822431e-37 = -4.9865316e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100100000000100101011001110100;
		b = 32'b11000011010111000100011000000011;
		correct = 32'b01100000000101110111101000110110;
		#400 //-9.617225e+21 * -220.27348 = 4.3660384e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000001100010110111011101010110;
		b = 32'b00111000001010010101100111111111;
		correct = 32'b00001000110100101101001011100100;
		#400 //5.1231775e-38 * 4.0376555e-05 = 1.2688495e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110101100001100001101111011011;
		b = 32'b01010111100111000000010100111111;
		correct = 32'b11011101010111000000110000001110;
		#400 //-3.4000623e+32 * 343092700000000.0 = -9.91004e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111000010010001100111000100111;
		b = 32'b01101110111111001111110001000101;
		correct = 32'b11001000110010110011001010110101;
		#400 //-1.629126e+34 * 3.9147599e+28 = -416149.66
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010111001001100010101101011110;
		b = 32'b10100110000011101010111001000000;
		correct = 32'b11110000100101010001001001101011;
		#400 //182705190000000.0 * -4.95023e-16 = -3.6908426e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010001010001000001110110011101;
		b = 32'b01001000101100011000111101101000;
		correct = 32'b10001000000011010110000001010111;
		#400 //-1.5470799e-28 * 363643.25 = -4.254389e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111001100100101000011011001000;
		b = 32'b01001110010110101000000010010010;
		correct = 32'b10101010101010111010110000011100;
		#400 //-0.0002794771 * 916464800.0 = -3.0495127e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000110010101111111111011111001;
		b = 32'b11011110110101100101101010101000;
		correct = 32'b10100111000000001111101011111101;
		#400 //13823.743 * -7.7229213e+18 = -1.789963e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101110110100001010111111111111;
		b = 32'b00010010101011001011000011101000;
		correct = 32'b01011011100110101010111001001101;
		#400 //9.490008e-11 * 1.0898337e-27 = 8.7077584e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100011100000110101001011110110;
		b = 32'b11010011001110100100111111101100;
		correct = 32'b10001111101101000111000110111001;
		#400 //1.4238184e-17 * -800204800000.0 = -1.7793175e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101010010110011101011011101111;
		b = 32'b00101100110111101000011011001010;
		correct = 32'b11111100111110101001101110101000;
		#400 //-6.5837975e+25 * 6.324584e-12 = -1.04098504e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111100100110011000110101010001;
		b = 32'b01111010101011111111011011111001;
		correct = 32'b11000001010111110110010010100101;
		#400 //-6.378301e+36 * 4.5683058e+35 = -13.962071
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011000100100001000010110101110;
		b = 32'b11101010100101100101110111101011;
		correct = 32'b10101101011101100000110010100110;
		#400 //1271230600000000.0 * -9.089119e+25 = -1.39862896e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111010111111100110001101101000;
		b = 32'b00010000011001011011001110000110;
		correct = 32'b01101010000011011100000110111010;
		#400 //0.0019408287 * 4.5300587e-29 = 4.2843347e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100110010110101111001011010111;
		b = 32'b01001101110101001001010000110010;
		correct = 32'b10011000000000111101010111011100;
		#400 //-7.5963053e-16 * 445810240.0 = -1.7039325e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101100001011001111101001000010;
		b = 32'b10111000110111100011000111011110;
		correct = 32'b10110010110001110100101101110101;
		#400 //2.4581591e-12 * -0.000105950734 = -2.3200963e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110001111011111011010100101010;
		b = 32'b01010110100011010110010110110001;
		correct = 32'b10011010110110001111111011100010;
		#400 //-6.9764114e-09 * 77733950000000.0 = -8.974729e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110010011011111110000100011011;
		b = 32'b11111010010000001111101101110010;
		correct = 32'b00110111100111110001101100001010;
		#400 //-4.7512994e+30 * -2.5050523e+35 = 1.8966868e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100001100110110000010111110110;
		b = 32'b11010000110101111000111010100111;
		correct = 32'b11010000001110000001101111010011;
		#400 //3.5745936e+20 * -28931602000.0 = -12355325000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111111000010110010011101100101;
		b = 32'b01110001010110001001111100111110;
		correct = 32'b10001101001001000111001100010101;
		#400 //-0.54356986 * 1.0726604e+30 = -5.0674927e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011111010010001100011010001011;
		b = 32'b11010110100000000111000110010101;
		correct = 32'b01001000010010000001010100000000;
		#400 //-1.4467404e+19 * -70612660000000.0 = 204884.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000101010110000001111001100001;
		b = 32'b00000101101101101011101101110110;
		correct = 32'b00111111000101110110001011101110;
		#400 //1.0161851e-35 * 1.718406e-35 = 0.5913533
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001101011000011101000111001000;
		b = 32'b00000101101011111011101110111110;
		correct = 32'b11000111001001000111101101000101;
		#400 //-6.9585993e-31 * 1.6525886e-35 = -42107.27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100001001000011010101111110001;
		b = 32'b10001001111010111010101011110010;
		correct = 32'b01010110101011111001111010110000;
		#400 //-5.4776484e-19 * -5.673495e-33 = 96548050000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100100101110110111001000010000;
		b = 32'b00010010110000001001101011011011;
		correct = 32'b11010001011110010010010001111001;
		#400 //-8.129155e-17 * 1.2155078e-27 = -66878673000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101111101111010010110100111101;
		b = 32'b01000111011001101101001001101110;
		correct = 32'b11100111110100011100111111100011;
		#400 //-1.1709471e+29 * 59090.43 = -1.9816189e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110101111011101100100001001011;
		b = 32'b10100001011101011010011110101001;
		correct = 32'b01010011111110001101011010001011;
		#400 //-1.7790675e-06 * -8.3231125e-19 = 2137502600000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101111001100100010000110000110;
		b = 32'b01100001010101110110000110010110;
		correct = 32'b10001101010100111011100110000111;
		#400 //-1.6200916e-10 * 2.4831761e+20 = -6.5242715e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001000000010101001101000101001;
		b = 32'b01010000010011100001010110100010;
		correct = 32'b00110111001011000010110001000001;
		#400 //141928.64 * 13830097000.0 = 1.0262303e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111001111110011100100101010010;
		b = 32'b11010101111100011011011011001100;
		correct = 32'b11100011100001000100011001010101;
		#400 //1.6212065e+35 * -33220926000000.0 = -4.8800763e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011100110110011110100010001;
		b = 32'b01001011100010000100110110010011;
		correct = 32'b10111111100100011100100000110100;
		#400 //-20347426.0 * 17865510.0 = -1.1389222
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001111000101110011101000111011;
		b = 32'b10110100000100110101011001001100;
		correct = 32'b00011010100000110110000100111001;
		#400 //-7.4560896e-30 * -1.3721836e-07 = 5.43374e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101100011011101111011010110100;
		b = 32'b01000001110100110100010000000111;
		correct = 32'b01101010000100001100100000001011;
		#400 //1.1555575e+27 * 26.408216 = 4.37575e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011001110000110011011001100011;
		b = 32'b00100000011001101001101010000110;
		correct = 32'b11111000110110001011011000010010;
		#400 //-6868427400000000.0 * 1.9532885e-19 = -3.5163405e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100001011100001010100110011100;
		b = 32'b10110111110001001111011001110101;
		correct = 32'b11101001000111000110011000101111;
		#400 //2.7746501e+20 * -2.3479786e-05 = -1.1817186e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011101000011011101010001101001;
		b = 32'b10101001010010011001010010101100;
		correct = 32'b10110011001101000001111001010010;
		#400 //1.8771008e-21 * -4.4759918e-14 = -4.1937092e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101010000010001100100011011000;
		b = 32'b01010100110001111000011100011100;
		correct = 32'b00010100101011110111111110100100;
		#400 //1.2148908e-13 * 6855722000000.0 = 1.772083e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101011110100011100000110110001;
		b = 32'b00011011011111011100000111011010;
		correct = 32'b01001111110100111001110001001001;
		#400 //1.4904103e-12 * 2.0990306e-22 = 7100470000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100101111000101100010110000010;
		b = 32'b10010101000100001111010010101101;
		correct = 32'b11010000010010000011111011100000;
		#400 //3.9338587e-16 * -2.9273584e-26 = -13438255000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000010111000000110001010000000;
		b = 32'b00100110110100111011100011011111;
		correct = 32'b00011011100001111010011111000111;
		#400 //3.2970378e-37 * 1.4691176e-15 = 2.24423e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010001111001111101100100111000;
		b = 32'b00111101100001000101111001100010;
		correct = 32'b00010011111000000011001001010101;
		#400 //3.6579245e-28 * 0.064633146 = 5.659518e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100011100100010001110110001;
		b = 32'b01010111110010111000000010000110;
		correct = 32'b00101100000110000100110101101001;
		#400 //968.5577 * 447505730000000.0 = 2.164347e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100110010101101011011110000100;
		b = 32'b01000011110100000000000111010100;
		correct = 32'b11100010000001000010000100000001;
		#400 //-2.5349292e+23 * 416.01428 = -6.093371e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101110001101000110100100100110;
		b = 32'b00111111000110111001100010111101;
		correct = 32'b11101110100101000110100110111111;
		#400 //-1.3958605e+28 * 0.60779935 = -2.296581e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010100010110111101101101101010;
		b = 32'b01111101010001111100000100110100;
		correct = 32'b10010110100011001110000110011111;
		#400 //-3777116000000.0 * 1.6594971e+37 = -2.2760607e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001110101000111000111111110110;
		b = 32'b10100111101010100001101010101001;
		correct = 32'b01100110011101100010011110100101;
		#400 //-1372060400.0 * -4.7213384e-15 = 2.9060837e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001111100101000100010010111110;
		b = 32'b01010101011010101011111101111100;
		correct = 32'b00111001101000011011000100000011;
		#400 //4975066000.0 * 16131759000000.0 = 0.00030840197
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001011010100000110000010001111;
		b = 32'b01001010011100100101000000000001;
		correct = 32'b01000000010111000010010111010100;
		#400 //13656207.0 * 3970048.2 = 3.4398088
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100011011100001010100111111010;
		b = 32'b11001010101001000111000110100000;
		correct = 32'b00011000001110110101010000001100;
		#400 //-1.304642e-17 * -5388496.0 = 2.4211616e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101110100101001100101000100010;
		b = 32'b10111011101000000000100011001001;
		correct = 32'b10110010011011100000001100100101;
		#400 //6.766167e-11 * -0.00488386 = -1.3854138e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100101110100100111101010000111;
		b = 32'b11000010111111010011110101101010;
		correct = 32'b01100010010101001100010111001101;
		#400 //-1.2424465e+23 * -126.61995 = 9.812407e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111100000110011100000101000110;
		b = 32'b11111000010011100001100111010100;
		correct = 32'b00000011001111101111101100001001;
		#400 //-0.009384459 * -1.6720891e+34 = 5.6124156e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000101101010110110011010101100;
		b = 32'b11000110001100111001010011000100;
		correct = 32'b00111110111101000101011011001001;
		#400 //-5484.834 * -11493.191 = 0.47722462
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010110101010010101111101011111;
		b = 32'b11000101100011011001100111010010;
		correct = 32'b11010000100110010001101010101100;
		#400 //93113540000000.0 * -4531.2275 = -20549296000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011000110100010000001010000000;
		b = 32'b11001111001111001000000100100101;
		correct = 32'b01001001000011011110110001110111;
		#400 //-1838469300000000.0 * -3162580200.0 = 581319.44
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000001001111110110001001100001;
		b = 32'b10011010010000011110110111100010;
		correct = 32'b10100110011111001010001111111000;
		#400 //3.5151743e-38 * -4.0103625e-23 = -8.765228e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010001110011010110001010101101;
		b = 32'b01011110111011000011110111110101;
		correct = 32'b10110010010111101001000000010001;
		#400 //-110265475000.0 * 8.511516e+18 = -1.2954858e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111111111000001010110100010110;
		b = 32'b00011111110000111110000111010110;
		correct = 32'b01011111100100101101000011000110;
		#400 //1.7552822 * 8.2959327e-20 = 2.1158346e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000001010001100100000101001010;
		b = 32'b10111001111001101111101100111110;
		correct = 32'b10000110110110111011101010011000;
		#400 //3.64137e-38 * -0.0004405621 = -8.265282e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000110001110110100100111111011;
		b = 32'b01011000111010101101000001110100;
		correct = 32'b10101100110011000010111111010100;
		#400 //-11986.495 * 2065448200000000.0 = -5.8033387e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001100011010100000000110101100;
		b = 32'b11011101100011110011001010100001;
		correct = 32'b10101110010100010010101111001110;
		#400 //61343410.0 * -1.2898108e+18 = -4.7560005e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110100000101001010101101010111;
		b = 32'b01000101000110011011101001111111;
		correct = 32'b10101110011101111001001100110110;
		#400 //-1.3845907e-07 * 2459.656 = -5.6292047e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010100101011110010011000000000;
		b = 32'b10010100111010101010011011101100;
		correct = 32'b11111111001111110001010100111011;
		#400 //6018054500000.0 * -2.3693801e-26 = -2.5399278e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010001101001011110101100010100;
		b = 32'b10001111011110011100111010001111;
		correct = 32'b01000001101010100000100000011011;
		#400 //-2.6177288e-28 * -1.23164296e-29 = 21.253958
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111000101111000111010100000101;
		b = 32'b01110100101110011110101110001001;
		correct = 32'b10000011100000011011111100100110;
		#400 //-8.986335e-05 * 1.1784084e+32 = -7.625824e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110011100101000011110101000010;
		b = 32'b01000111110110000100011111101100;
		correct = 32'b10101011001011110111011001111001;
		#400 //-6.90293e-08 * 110735.84 = -6.2336903e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011110001001110000010110011;
		b = 32'b10100010010000011001110101110011;
		correct = 32'b01101001000000100010100000110000;
		#400 //-25805158.0 * -2.623973e-18 = 9.834384e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101101010100010111110100001101;
		b = 32'b01100101010001100000001001111100;
		correct = 32'b10000111100001110110101110010110;
		#400 //-1.1908041e-11 * 5.844215e+22 = -2.0375776e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010101111100100001111100110011;
		b = 32'b10011100100101000101011100100101;
		correct = 32'b00111000110100001110110000010011;
		#400 //-9.7792245e-26 * -9.816345e-22 = 9.962185e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000011111010001100101001000111;
		b = 32'b11101000110010110101100001001110;
		correct = 32'b10011010100100101000100011110010;
		#400 //465.5803 * -7.6821546e+24 = -6.060543e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010010110110100001011111100000;
		b = 32'b11111000111000100010100111111011;
		correct = 32'b00011001011101101101110101010100;
		#400 //-468351700000.0 * -3.6697205e+34 = 1.2762599e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111101010111111111110110100000;
		b = 32'b11001010101111111010101000011001;
		correct = 32'b11110010000101011001011010101101;
		#400 //1.8608421e+37 * -6280460.5 = -2.962907e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100100100011101110100110100011;
		b = 32'b11000000010010001010010010100010;
		correct = 32'b01100011101101100101011110000101;
		#400 //-2.1090184e+22 * -3.1350484 = 6.727228e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100100010010111001101100110010;
		b = 32'b00000011010001001110000001100101;
		correct = 32'b01100000100001000110000000010110;
		#400 //4.4150064e-17 * 5.7856815e-37 = 7.6309186e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110010001111110011010101111000;
		b = 32'b11010011101001110100011000001011;
		correct = 32'b00011110000100100101000011001010;
		#400 //-1.1129821e-08 * -1436869300000.0 = 7.7458824e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010110100010010111111000100100;
		b = 32'b11001011111011001101100011110000;
		correct = 32'b01001010000101001001110001101101;
		#400 //-75587430000000.0 * -31044064.0 = 2434843.2
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101101110100100110001010000011;
		b = 32'b00111000100001000110010011100001;
		correct = 32'b10110100110010110110011011111101;
		#400 //-2.3917984e-11 * 6.313041e-05 = -3.788663e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100001101001110011111001101101;
		b = 32'b00100000010111001011011111010001;
		correct = 32'b01000000110000011111101001011001;
		#400 //1.1332884e-18 * 1.8695545e-19 = 6.06181
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101011001110111000000101000101;
		b = 32'b10110000010111111110110001100101;
		correct = 32'b11111010010101100101110101011011;
		#400 //2.2667959e+26 * -8.1462864e-10 = -2.7826125e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111100010000001101011010101101;
		b = 32'b01100001001011100111010010101101;
		correct = 32'b00011010100011010111110011010111;
		#400 //0.011769933 * 2.011338e+20 = 5.851792e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011001010100001000000100101000;
		b = 32'b11001111100010110010110010111110;
		correct = 32'b11001001001111111100001101010111;
		#400 //3668050200000000.0 * -4669930500.0 = -785461.44
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001011110111101000010010100101;
		b = 32'b00001010110010100110000110010101;
		correct = 32'b11000000100011001011110001101100;
		#400 //-8.571087e-32 * 1.9488599e-32 = -4.3980007
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001011010000000101110111110111;
		b = 32'b00001001000100100110010101110010;
		correct = 32'b11000001101010000011000110101110;
		#400 //-3.7048546e-32 * 1.762181e-33 = -21.024258
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000111101100000000011111010110;
		b = 32'b11011000110111111101100000010111;
		correct = 32'b00101110010010010101000101100101;
		#400 //-90127.67 * -1968953500000000.0 = 4.57744e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100100011100010010010010001111;
		b = 32'b00111001011110011111110011000110;
		correct = 32'b01101010011101101111000101010100;
		#400 //1.7793199e+22 * 0.00023840656 = 7.463385e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000100101111100111000111011110;
		b = 32'b10000001100000100001100011000001;
		correct = 32'b01000010101110110110000000100001;
		#400 //-4.4773356e-36 * -4.778998e-38 = 93.68775
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100011011001001010101000101100;
		b = 32'b11000110101110011010111000000001;
		correct = 32'b01011100000111011010000111010011;
		#400 //-4.2181198e+21 * -23767.002 = 1.77478e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100011000011001010010011010011;
		b = 32'b01101010001110000101111110010010;
		correct = 32'b10111000010000110100100000111101;
		#400 //-2.594421e+21 * 5.5723417e+25 = -4.65589e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000000011100010001111110111011;
		b = 32'b11110100111001111100111111011010;
		correct = 32'b00001011000001010010010001010000;
		#400 //-3.7675617 * -1.4692826e+32 = 2.5642187e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101100011010001001010010011110;
		b = 32'b11111110011010100101100011111011;
		correct = 32'b00101101011111100001000111010111;
		#400 //-1.12469046e+27 * -7.787534e+37 = 1.444219e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101011011100010110101001011001;
		b = 32'b01001001100100011011011110101001;
		correct = 32'b10100001010101000000111111110100;
		#400 //-8.5767987e-13 * 1193717.1 = -7.184951e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000100100100000101010110110;
		b = 32'b10101000011100100111010010111101;
		correct = 32'b01000111100110100011001100110010;
		#400 //-1.0625942e-09 * -1.3459012e-14 = 78950.39
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100011111011100111110011101110;
		b = 32'b01001011001101010011010011111011;
		correct = 32'b01011000001010000111011000111110;
		#400 //8.7986544e+21 * 11875579.0 = 740903200000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110011100010011101011110101110;
		b = 32'b10011101111001110010111001111010;
		correct = 32'b01010101000110001010001111111011;
		#400 //-6.4187915e-08 * -6.1193247e-21 = 10489379000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001110100110100110000111100101;
		b = 32'b00010101110010110111111010100111;
		correct = 32'b00111000010000100011011100111111;
		#400 //3.80582e-30 * 8.219087e-26 = 4.6304656e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111101000100010111010010010001;
		b = 32'b11001001010101011100101110100101;
		correct = 32'b01110011001011100010101101001010;
		#400 //-1.2083957e+37 * -875706.3 = 1.3799098e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001100000110010101100110011100;
		b = 32'b00110111110100000100110111000100;
		correct = 32'b01010011101111000111011010011001;
		#400 //40199790.0 * 2.4831745e-05 = 1618887200000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101011000101101011101110101110;
		b = 32'b10010110011111001111110101001111;
		correct = 32'b01010100000110001000011011011101;
		#400 //-5.3551163e-13 * -2.0436328e-25 = 2620390600000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001111110000001011110111110010;
		b = 32'b00010100011001000001110001100111;
		correct = 32'b11111010110110000100111010001001;
		#400 //-6467347500.0 * 1.151666e-26 = -5.615645e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001001000001001110010100111001;
		b = 32'b01101000110110111010101110110011;
		correct = 32'b10011111100110101101111110101101;
		#400 //-544339.56 * 8.2989244e+24 = -6.559158e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001011111101011011101111101000;
		b = 32'b10111100011100011100010111101001;
		correct = 32'b00001111000000100001100011010101;
		#400 //-9.46533e-32 * -0.014756658 = 6.414277e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110001101111111100101110110101;
		b = 32'b00101110010111001100010111001001;
		correct = 32'b01000010110111100110011001000011;
		#400 //5.5819904e-09 * 5.0197877e-11 = 111.19973
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101001000001111101110011110011;
		b = 32'b00001000000010011001000110101111;
		correct = 32'b11100000011111001101001101001010;
		#400 //-3.0167665e-14 * 4.139819e-34 = -7.2871945e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110101001011011011101111110001;
		b = 32'b01110010000001001001100101000111;
		correct = 32'b10000010101001111011010101110010;
		#400 //-6.4721013e-07 * 2.6263886e+30 = -2.464259e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010001101101111000101111011100;
		b = 32'b11100001011111100011001001110000;
		correct = 32'b10101111101110001101100100100011;
		#400 //98540680000.0 * -2.9306921e+20 = -3.362369e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001011101011110010100001000000;
		b = 32'b11001101101101100111110011010101;
		correct = 32'b10111101011101011011011101110111;
		#400 //22958208.0 * -382704300.0 = -0.05998942
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011101010001011111010010110000;
		b = 32'b01100110100010010010110000100111;
		correct = 32'b00110110001110001011100000001000;
		#400 //8.915137e+17 * 3.2388934e+23 = 2.7525257e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110010001101111100110111111101;
		b = 32'b01000110100101001000000111100100;
		correct = 32'b11101011000111100110110001001110;
		#400 //-3.640626e+30 * 19008.945 = -1.9152173e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100101000101110110100010010110;
		b = 32'b10011010110011101000111011000011;
		correct = 32'b11001001101110111010011001110011;
		#400 //1.3132597e-16 * -8.543025e-23 = -1537230.4
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000001110000111011000011101110;
		b = 32'b00011010011011010111000110010111;
		correct = 32'b10100110110100101111110000000101;
		#400 //-7.188557e-38 * 4.910221e-23 = -1.4639987e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000100101110100010111100010111;
		b = 32'b10001110011100001100010111011000;
		correct = 32'b01110101110001011111010101110001;
		#400 //-1489.4716 * -2.9677542e-30 = 5.0188507e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111011010111111111000001111111;
		b = 32'b01110101001111001111101110110010;
		correct = 32'b00000101100101111010110100011010;
		#400 //0.0034170446 * 2.3956465e+32 = 1.4263559e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101101100111101101110011000010;
		b = 32'b10111011010101001110101100111100;
		correct = 32'b10110001101111110000000110000001;
		#400 //1.8060557e-11 * -0.0032488843 = -5.5590026e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100001010000010101011100110001;
		b = 32'b11010111000010001110110010110101;
		correct = 32'b11001001101101001011110100100011;
		#400 //2.2290653e+20 * -150550230000000.0 = -1480612.4
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011011100010110011101110011111;
		b = 32'b11011000001101110001100000111111;
		correct = 32'b01000010110000101010110001010010;
		#400 //-7.838115e+16 * -805259060000000.0 = 97.33656
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110100110101100011011000011101;
		b = 32'b00000011111000010001100101100111;
		correct = 32'b11110000011100111001111000010101;
		#400 //-3.989998e-07 * 1.32301435e-36 = -3.0158387e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011001011101110110111110111101;
		b = 32'b00101011111101110101101011011111;
		correct = 32'b01101101000000000000101011001100;
		#400 //4352948500000000.0 * 1.7575627e-12 = 2.476696e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101111000101010100001101101001;
		b = 32'b10101000001010100011100101010111;
		correct = 32'b11000110011000000111101000101100;
		#400 //1.357542e-10 * -9.449329e-15 = -14366.543
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011011010101100100101010101;
		b = 32'b00011111011010100011110011101001;
		correct = 32'b11101011100000000100110010111100;
		#400 //-15386965.0 * 4.960181e-20 = -3.1020975e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110010010111000010101100000110;
		b = 32'b01111001101001111111111111000111;
		correct = 32'b00111000001001111011111101111010;
		#400 //4.3608777e+30 * 1.0903767e+35 = 3.999423e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011110011100011011010011010111;
		b = 32'b11001011101011010010010010011101;
		correct = 32'b01010010001100101010111111100100;
		#400 //-4.3541955e+18 * -22694202.0 = 191863780000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111010100011001100100111011110;
		b = 32'b11100100100111110100000111010100;
		correct = 32'b01010101011000100100111111111010;
		#400 //-3.6550796e+35 * -2.3502206e+22 = 15552070000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011111000101110011010011111000;
		b = 32'b00111101101100111011010001001011;
		correct = 32'b10100000110101110110011101011010;
		#400 //-3.201931e-20 * 0.087746225 = -3.649081e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010011110110010110100011111111;
		b = 32'b10101011000011011100010110111001;
		correct = 32'b00101000010001000100101000111111;
		#400 //-5.4882035e-27 * -5.036766e-13 = 1.0896285e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010110010110011000110011000110;
		b = 32'b11100100000100101110100010010111;
		correct = 32'b10110001101111011000110010010011;
		#400 //59799660000000.0 * -1.0839938e+22 = -5.5166054e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010100000111000011000111010000;
		b = 32'b11001011111100001001111001101111;
		correct = 32'b10000111101001100010110111010101;
		#400 //7.885811e-27 * -31538398.0 = -2.5003842e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111010000100100100110000101101;
		b = 32'b01000001000000001111111010011011;
		correct = 32'b11111000100100010010101101101011;
		#400 //-1.899051e+35 * 8.06216 = -2.3555115e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011100110000011000100011011000;
		b = 32'b11000110010011101001110000011001;
		correct = 32'b00010101111011111100110010010101;
		#400 //-1.2807042e-21 * -13223.024 = 9.6854105e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000101100111010001111110101101;
		b = 32'b01110001000000110101111110000111;
		correct = 32'b10010100000110010001011011100011;
		#400 //-5027.9595 * 6.5052835e+29 = -7.7290396e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100011000100011001111101000110;
		b = 32'b00001001000100100000000000111100;
		correct = 32'b01011001011111110101010111111101;
		#400 //7.894193e-18 * 1.7574221e-33 = 4491916500000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101110011101111011111101110011;
		b = 32'b10010110001110010101010100010100;
		correct = 32'b01010111101010110001101101111011;
		#400 //-5.633134e-11 * -1.4971027e-25 = 376269030000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101001011110101011100100011100;
		b = 32'b10000101101010110100010001011000;
		correct = 32'b11100011001110110110001000011010;
		#400 //5.5671708e-14 * -1.6105868e-35 = -3.45661e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010110010001100001111110101000;
		b = 32'b00100011101011001000000001101100;
		correct = 32'b00110010000100110000001100011000;
		#400 //1.6004302e-25 * 1.8702666e-17 = 8.55723e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010110001001000011010010010101;
		b = 32'b01001000111011110110000010101000;
		correct = 32'b10001100101011111001101110011101;
		#400 //-1.3264406e-25 * 490245.25 = -2.7056676e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001101010010110011101111111101;
		b = 32'b11010100011111010100010101011000;
		correct = 32'b10111000010011010110110010011110;
		#400 //213106640.0 * -4351160500000.0 = -4.8976966e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001000011000001110110010101110;
		b = 32'b00001101100000000010111110010110;
		correct = 32'b10111010011000001001100100101111;
		#400 //-6.7685764e-34 * 7.900065e-31 = -0.0008567748
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010100111010010110001101010100;
		b = 32'b01001110000100100100010100110010;
		correct = 32'b10000110010011000011110001101100;
		#400 //-2.3566166e-26 * 613502100.0 = -3.8412527e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111111111100111001101101001010;
		b = 32'b11011001011111101110111101101110;
		correct = 32'b01111111111100111001101101001010;
		#400 //nan * -4484868700000000.0 = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110111111001011000000101011111;
		b = 32'b11100101010111101000010001001011;
		correct = 32'b01010010000001000000010100100101;
		#400 //-9.309843e+33 * -6.567536e+22 = 141755500000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011111110111010100010110111011;
		b = 32'b10111001000011101101011001111001;
		correct = 32'b11100110010001100100100101110100;
		#400 //3.1888711e+19 * -0.00013622073 = -2.3409588e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000110100011101111000000101001;
		b = 32'b00100110000110111111001001100111;
		correct = 32'b01011111111010101010010100100000;
		#400 //18296.08 * 5.4104944e-16 = 3.3815911e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100110001111011111110100011111;
		b = 32'b11000101001110010000100001111100;
		correct = 32'b10100000100000110110110110011010;
		#400 //6.591559e-16 * -2960.5303 = -2.2264791e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100110011000001101100011101111;
		b = 32'b10001011110110100110100010111100;
		correct = 32'b11011010000000111100010111110000;
		#400 //7.800961e-16 * -8.412813e-32 = -9272714000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101101101010001110010110100010;
		b = 32'b01111100101011111010010110101001;
		correct = 32'b10110000011101100010100101110101;
		#400 //-6.5338863e+27 * 7.2960955e+36 = -8.955319e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100111111010011111110110000000;
		b = 32'b01001111110110010110100111001011;
		correct = 32'b10010111100010011100001001110001;
		#400 //-6.4945336e-15 * 7295178000.0 = -8.902501e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011110101101111000001000001101;
		b = 32'b00111111010100000011100111111100;
		correct = 32'b11011110111000011001110000111111;
		#400 //-6.611573e+18 * 0.8133848 = -8.128469e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101000000111101011100111101001;
		b = 32'b01001000001000010101010011100100;
		correct = 32'b11011111011110111101110110100100;
		#400 //-2.9982534e+24 * 165203.56 = -1.8148842e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111001001110100111111101001000;
		b = 32'b11111110010000001110010101111010;
		correct = 32'b10111010011101111000000111100100;
		#400 //6.05218e+34 * -6.410082e+37 = -0.00094416575
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101010101111100111001000110011;
		b = 32'b00010001011011110111010111010110;
		correct = 32'b11011000110010111001100110110000;
		#400 //-3.3830022e-13 * 1.8890087e-28 = -1790887500000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100111000110010101101100110001;
		b = 32'b00111111111001101010100101001101;
		correct = 32'b00100110101010100011001111100111;
		#400 //2.128245e-15 * 1.8020416 = 1.1810188e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000100110111101111010010000000;
		b = 32'b10001111100110010111111011101000;
		correct = 32'b00110100101110011110110000010000;
		#400 //-5.2416487e-36 * -1.5135847e-29 = 3.4630693e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111110001011000010111110110011;
		b = 32'b10011111110101001010110010001111;
		correct = 32'b01011101110011110100001110011101;
		#400 //-0.16815071 * -9.0070967e-20 = 1.8668692e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111001010001100110010000101011;
		b = 32'b01010000000011001101011100101100;
		correct = 32'b00101000101101000100110111001000;
		#400 //0.00018920067 * 9451647000.0 = 2.0017747e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010100011000010101000001011110;
		b = 32'b00101010011011000010111110010011;
		correct = 32'b11101001011101000011011101001110;
		#400 //-3870864000000.0 * 2.0977516e-13 = -1.8452442e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011010111000011101001101110101;
		b = 32'b10000110001000000100010100100010;
		correct = 32'b11010100001101000101101100111101;
		#400 //9.3399446e-23 * -3.0143446e-35 = -3098499400000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111111101111011110110111010110;
		b = 32'b00001100001110101011110000101000;
		correct = 32'b01110011000000100011000001111101;
		#400 //1.4838207 * 1.438554e-31 = 1.0314668e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000001110101101111010010100100;
		b = 32'b01110011011100001000010001100011;
		correct = 32'b10001101111001001100101100000011;
		#400 //-26.869453 * 1.9055731e+31 = -1.4100458e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000001000010010000110001111101;
		b = 32'b00010110101010111110100011001101;
		correct = 32'b01101001110011000001011001001101;
		#400 //8.565549 * 2.7773458e-25 = 3.0840772e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111001111000101011110101001011;
		b = 32'b01011010110010101111110101010100;
		correct = 32'b11011110100011101111100111011111;
		#400 //-1.471623e+35 * 2.8568241e+16 = -5.1512554e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100001111011001010011000011010;
		b = 32'b01000111101001000100001000011000;
		correct = 32'b00011001101110000110100101000110;
		#400 //1.6035949e-18 * 84100.19 = 1.9067674e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000101001101110101011100001101;
		b = 32'b11110010101110100100111101001101;
		correct = 32'b10010001111110111110101101100000;
		#400 //2933.4407 * -7.3804903e+30 = -3.9745878e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010100011101100100010111111001;
		b = 32'b10100101101011111101000101111110;
		correct = 32'b11101110001100110100101011111111;
		#400 //4230943600000.0 * -3.0499618e-16 = -1.387212e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110100001011100010011011000011;
		b = 32'b01011001011101000110100100001101;
		correct = 32'b01011010001101100110100011010011;
		#400 //5.5190786e+31 * 4299712400000000.0 = 1.2835925e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100000001110110100111101111100;
		b = 32'b00011001001110000110001011001001;
		correct = 32'b01000110100000100000011110111111;
		#400 //1.5865815e-19 * 9.5325265e-24 = 16643.873
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011000011101001000000010011010;
		b = 32'b11011110110100010100011001101011;
		correct = 32'b00111001000101011000101111010111;
		#400 //-1075332700000000.0 * -7.539929e+18 = 0.00014261842
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110001011000000101111001000010;
		b = 32'b10010101100000001100000110001011;
		correct = 32'b11011011010111110000110011111110;
		#400 //3.264987e-09 * -5.2004145e-26 = -6.2783205e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101010011111110010011000011101;
		b = 32'b01100001110010100001100000110010;
		correct = 32'b10001000001000011001101001010111;
		#400 //-2.2661773e-13 * 4.6599822e+20 = -4.86306e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111101011000000111111011010111;
		b = 32'b11100000011001101101010011000100;
		correct = 32'b11011100011110001111100100111010;
		#400 //1.8650354e+37 * -6.653254e+19 = -2.8031929e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010111110111101101010011101100;
		b = 32'b01001101011101010000110111110000;
		correct = 32'b01001001111010001100100011100001;
		#400 //490012150000000.0 * 256958200.0 = 1906972.1
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100010100100101101001001010000;
		b = 32'b00110101001101000001000000111010;
		correct = 32'b11101100110100001011110101000110;
		#400 //-1.3541896e+21 * 6.707884e-07 = -2.0188031e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000001011100000011011111000101;
		b = 32'b00111101100100000010110101100100;
		correct = 32'b01000011010101010100001110101111;
		#400 //15.013616 * 0.070399076 = 213.26439
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111000001000100101100011110101;
		b = 32'b11011100110110100100110010001101;
		correct = 32'b10011010101111100110001010101100;
		#400 //3.8706658e-05 * -4.915657e+17 = -7.874157e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100011110001001111000110101111;
		b = 32'b10110011111111111010101101001011;
		correct = 32'b00101111010001010011001011101111;
		#400 //-2.135272e-17 * -1.1905521e-07 = 1.7935141e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100001101011110100000101001010;
		b = 32'b00011110100010011001000000010011;
		correct = 32'b11000010101000110001001001110001;
		#400 //-1.1875743e-18 * 1.4565027e-20 = -81.53602
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101111100101001101100000011100;
		b = 32'b00010001111001101110011010111110;
		correct = 32'b11011101001001010000010111111001;
		#400 //-2.7074598e-10 * 3.6429807e-28 = -7.43199e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011111001000001111000101011111;
		b = 32'b10001001100100011000001100010001;
		correct = 32'b11010101000011011001001011100101;
		#400 //3.4080975e-20 * -3.5030734e-33 = -9728878000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000010100010100001110111110;
		b = 32'b11001000100000010110101100001000;
		correct = 32'b00100111010011101111100010111100;
		#400 //-7.6130025e-10 * -265048.25 = 2.8723082e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010101010001010010000100111111;
		b = 32'b00100010101000110111101110111011;
		correct = 32'b01110010000110100101011111111110;
		#400 //13546661000000.0 * 4.4312243e-18 = 3.0570923e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001100001010101110001000100111;
		b = 32'b01011000000011110011110110100010;
		correct = 32'b00110011100110001011001110010101;
		#400 //44796060.0 * 629979500000000.0 = 7.110717e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010111010001100010000111010110;
		b = 32'b01111101111010111001010101100000;
		correct = 32'b10011000110101110100110110010010;
		#400 //-217848630000000.0 * 3.9143022e+37 = -5.5654523e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100000001110111000001100000100;
		b = 32'b01001010111010110000000010010010;
		correct = 32'b01010100110011000100010000100111;
		#400 //5.404659e+19 * 7700553.0 = 7018534000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010011000010010011001001111001;
		b = 32'b10110011001100100010010110011001;
		correct = 32'b00011111010001010010011110010011;
		#400 //-1.7316716e-27 * -4.147805e-08 = 4.1749108e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000000010011101101011101010001;
		b = 32'b00110000100100010100011010100110;
		correct = 32'b01001111001101100011111001110000;
		#400 //3.2318919 * 1.0570218e-09 = 3057545200.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000101001101100110101001100000;
		b = 32'b00100011010000000010111111011101;
		correct = 32'b00100001011100101111101111101101;
		#400 //8.577137e-36 * 1.0418476e-17 = 8.232621e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001000110111001101011011000110;
		b = 32'b11111011100010100011001011100110;
		correct = 32'b00001100110011001000101010011100;
		#400 //-452278.2 * -1.4351386e+36 = 3.15146e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100010010010100110011001101101;
		b = 32'b10100101010101101100010101000011;
		correct = 32'b00111100011100010100000100111010;
		#400 //-2.7430329e-18 * -1.8628376e-16 = 0.014725024
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110001101010111001111111111011;
		b = 32'b10100011100011011101101101110101;
		correct = 32'b01001101100110101101110000011110;
		#400 //-4.9949427e-09 * -1.5380194e-17 = 324764600.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101010001101001110100011100101;
		b = 32'b00101101010000000101011110101010;
		correct = 32'b00111100011100001100100010010111;
		#400 //1.6068013e-13 * 1.0933402e-11 = 0.014696262
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111000100111110111010101000000;
		b = 32'b11011000100001001001101010001101;
		correct = 32'b01011111100110011110110000000110;
		#400 //-2.587354e+34 * -1166394600000000.0 = 2.2182493e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000000101111010100101110101;
		b = 32'b11000101000010010110100011101000;
		correct = 32'b00101010100011010100011010110011;
		#400 //-5.5174293e-10 * -2198.5566 = 2.509569e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010010011011000000111000000101;
		b = 32'b10110011111100001011110000101001;
		correct = 32'b01011101111110110000010111100011;
		#400 //-253461870000.0 * -1.1210097e-07 = 2.2610141e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001001101011101000011111101110;
		b = 32'b10011000100001100000000101000010;
		correct = 32'b00110000101001101011010111000101;
		#400 //-4.2016804e-33 * -3.463946e-24 = 1.2129752e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111111001101110001110111011000;
		b = 32'b00010011101000001110001110101001;
		correct = 32'b11101011000100011010111011111100;
		#400 //-0.7152991 * 4.061417e-27 = -1.7612058e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001001011111010100011010111000;
		b = 32'b11010101110001010001010111111001;
		correct = 32'b10110011001001000111111001011101;
		#400 //1037419.5 * -27087270000000.0 = -3.8299152e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000110000110011001001011000110;
		b = 32'b01000000100110111010110100011001;
		correct = 32'b11000100111111001000101011000010;
		#400 //-9828.693 * 4.86488 = -2020.3362
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000111011100111001000011000100;
		b = 32'b00100000001001111110110001010111;
		correct = 32'b11100110101110011010100010011000;
		#400 //-62352.766 * 1.4223649e-19 = -4.383739e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111010000000001010100111110001;
		b = 32'b00000000011111001010110000110000;
		correct = 32'b01111001000001000001100100000110;
		#400 //0.0004908136 * 1.1449371e-38 = 4.286817e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100111011000001010001110000000;
		b = 32'b10111110101110101000100011011001;
		correct = 32'b11101000000110100010010110100100;
		#400 //1.0608261e+24 * -0.3643253 = -2.911755e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110000100011001001000100010011;
		b = 32'b00110110000001000110101000100110;
		correct = 32'b11111010000001111110000101011001;
		#400 //-3.480263e+29 * 1.973132e-06 = -1.7638267e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100101000100010100111000111;
		b = 32'b01101111111010011000000000111000;
		correct = 32'b00010100001100011100100111011110;
		#400 //1297.3055 * 1.4453003e+29 = 8.976028e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111001110111010111001001111001;
		b = 32'b11110000101111100100011011000100;
		correct = 32'b01001000100101001111011111111110;
		#400 //-1.4372742e+35 * -4.711016e+29 = 305087.94
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101100111101000011001001101001;
		b = 32'b11110000010100100110011111001011;
		correct = 32'b00111100000101001000111010011001;
		#400 //-2.3617276e+27 * -2.6046932e+29 = 0.009067201
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111101101110100101011010011111;
		b = 32'b00011101001110000101001001101011;
		correct = 32'b11100000000000010110011001111000;
		#400 //-0.09098553 * 2.4394806e-21 = -3.729709e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001110110011100111011100110001;
		b = 32'b11001101010111110010010110100001;
		correct = 32'b11000000111011001101110011011000;
		#400 //1731958900.0 * -233986580.0 = -7.4019585
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101001100000100000011111110011;
		b = 32'b01001100000011011011111111111111;
		correct = 32'b10011100111010101101010111101101;
		#400 //-5.774539e-14 * 37158908.0 = -1.554012e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111111001110010110110010000011;
		b = 32'b11001011110111111101111110011100;
		correct = 32'b10110010110101000000100001100011;
		#400 //0.724312 * -29343544.0 = -2.4683862e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000110101111000011100101111;
		b = 32'b10001100111111011010001100011110;
		correct = 32'b01100011010110011000100100101111;
		#400 //-1.568173e-09 * -3.9078995e-31 = 4.0128286e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001110111110111110010011011110;
		b = 32'b01111110001000110011001010010101;
		correct = 32'b00010000010001011001000100011101;
		#400 //2113040100.0 * 5.42317e+37 = 3.896319e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001001010101001100101011101100;
		b = 32'b11111111000001111101110001010111;
		correct = 32'b10001001110010000111101100010101;
		#400 //871598.75 * -1.8058985e+38 = -4.8263994e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000010101010000110011000010101;
		b = 32'b11111110110110001111010011011010;
		correct = 32'b00000011010001101011010000101111;
		#400 //-84.19938 * -1.4419229e+38 = 5.839381e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111001001010010100110011011101;
		b = 32'b11011100100010000001000100111101;
		correct = 32'b11011100000111110100001100110111;
		#400 //5.494107e+34 * -3.063964e+17 = -1.793137e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110000110100100101101011100001;
		b = 32'b11001010010000101001000000000111;
		correct = 32'b10100110000010100110001110111100;
		#400 //1.530534e-09 * -3187713.8 = -4.8013533e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110011100110101110010100101010;
		b = 32'b00111001011100000101010010101110;
		correct = 32'b01111001101001001111111001111110;
		#400 //2.454412e+31 * 0.00022919729 = 1.070873e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110110101000010110011010101101;
		b = 32'b11011100001100101011011111111000;
		correct = 32'b01011001111001110011000110101010;
		#400 //-1.6368014e+33 * -2.0121929e+17 = 8134415700000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111101001000001000111010000001;
		b = 32'b11001010111010010011010101111011;
		correct = 32'b11110001101100000011111101100001;
		#400 //1.3338525e+37 * -7641789.5 = -1.7454714e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111010010001011100100010001010;
		b = 32'b01011111000100010010100000001011;
		correct = 32'b11011010101011100110100000100101;
		#400 //-2.5673747e+35 * 1.0459622e+19 = -2.4545577e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100011100101100100100010100101;
		b = 32'b10110110001010100111111001111011;
		correct = 32'b10101100111000011010011101100100;
		#400 //1.6293799e-17 * -2.5405595e-06 = -6.4134687e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000110110001101111010100011110;
		b = 32'b01000010011000000110001100110000;
		correct = 32'b11000011111000101111110011000100;
		#400 //-25466.559 * 56.096863 = -453.97473
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000101111110110101101101010011;
		b = 32'b01000111000011010001111000110101;
		correct = 32'b00111110011000111111110111000000;
		#400 //8043.4155 * 36126.207 = 0.22264767
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010100010010111011000111001001;
		b = 32'b00110111110100011101010000111101;
		correct = 32'b00011011111110001000001111111100;
		#400 //1.0283943e-26 * 2.5013573e-05 = 4.1113451e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001100100111000110000101001010;
		b = 32'b10011010100010111100101010010100;
		correct = 32'b11110001100011110011000010000001;
		#400 //81988180.0 * -5.7816335e-23 = -1.4180798e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111100101100000001011001111000;
		b = 32'b11011010101110100110100001000111;
		correct = 32'b10100001011100011101001111101000;
		#400 //0.021495089 * -2.62345e+16 = -8.193443e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011000100001011111000101101011;
		b = 32'b00001001001001001110101110101110;
		correct = 32'b01001110110011111110101000101000;
		#400 //3.4623464e-24 * 1.9851598e-33 = 1744114700.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010110001100111011010001010101;
		b = 32'b10100101111101000100101001000001;
		correct = 32'b11101111101111000101000110001000;
		#400 //49396775000000.0 * -4.237757e-16 = -1.1656349e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110011010111101110100001100111;
		b = 32'b01011001110001100100100011010111;
		correct = 32'b01011001000011111110010100101111;
		#400 //1.7660577e+31 * 6976516700000000.0 = 2531432000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010000010101101001101000110111;
		b = 32'b10100111011010111111010110110100;
		correct = 32'b00101000011010001101010000100111;
		#400 //-4.232286e-29 * -3.2745997e-15 = 1.292459e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010010111011100010100000000101;
		b = 32'b10010001000101110001100001011000;
		correct = 32'b11000001010010011100000011111001;
		#400 //1.5029777e-27 * -1.1919301e-28 = -12.609612
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111010101000100111011000101110;
		b = 32'b01001110111010111111011001110011;
		correct = 32'b11101011001100000100000111100111;
		#400 //-4.2177453e+35 * 1979398500.0 = -2.1308216e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010001110000010101100001100011;
		b = 32'b00010000110100000011011111010000;
		correct = 32'b01000000011011011011011011011000;
		#400 //3.0504503e-28 * 8.2127527e-29 = 3.714285
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011111010011111110110010010110;
		b = 32'b00010110111001101010101110111111;
		correct = 32'b01000111111001101100000101101100;
		#400 //4.4029654e-20 * 3.726689e-25 = 118146.84
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100001010011101000111101100100;
		b = 32'b10111011101110011001011010001101;
		correct = 32'b10100101000011100111011011100011;
		#400 //6.998529e-19 * -0.005663699 = -1.2356817e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110100100000110101001010110001;
		b = 32'b01110000110111111001110011011010;
		correct = 32'b01000011000101100101011111101000;
		#400 //8.323585e+31 * 5.5363823e+29 = 150.34338
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101000011100110011000110110011;
		b = 32'b10110000101001011000100110010001;
		correct = 32'b10110111001111000000110000011010;
		#400 //1.34999865e-14 * -1.2044429e-09 = -1.1208491e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111100110000111110111100111110;
		b = 32'b11000001011011111110110110110010;
		correct = 32'b01111010110100010000111100100011;
		#400 //-8.1388024e+36 * -14.995531 = 5.4274853e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011111100010000101100000000001;
		b = 32'b00101100010100000110111111111110;
		correct = 32'b11110010101001110111010010011101;
		#400 //-1.9649207e+19 * 2.9620746e-12 = -6.6335966e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011111001010100110001001110110;
		b = 32'b11111110000000101010000000101011;
		correct = 32'b00100000101001101111010110110100;
		#400 //-1.2277505e+19 * -4.340782e+37 = 2.8284087e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101110100000001011111110001010;
		b = 32'b00111001101011011000111010110111;
		correct = 32'b11110100001111011110011111010110;
		#400 //-1.992282e+28 * 0.00033103462 = -6.018349e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111010100000110011111000101110;
		b = 32'b01000100011111000011101011100100;
		correct = 32'b11110101100001010011010001011011;
		#400 //-3.4072602e+35 * 1008.92017 = -3.3771356e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111111101010000001010010110111;
		b = 32'b01000011000101011010101110011110;
		correct = 32'b00111100000011111011111010110011;
		#400 //1.3131322 * 149.67038 = 0.008773494
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000111001101101001101011011010;
		b = 32'b10001000100101000010000100101111;
		correct = 32'b00111110000111011100101001010101;
		#400 //-1.3737665e-34 * -8.915227e-34 = 0.15409215
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000000101001011000001110010;
		b = 32'b01101100100110111111101011110011;
		correct = 32'b10000010111101000000100010100010;
		#400 //-5.409283e-10 * 1.5085486e+27 = -3.5857533e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101001101011001110111101101000;
		b = 32'b10010010011010001001000001101110;
		correct = 32'b01010110101111100101110010110011;
		#400 //-7.679865e-14 * -7.3384315e-28 = 104652675000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101101000011111010011100010001;
		b = 32'b01111001001100101101110110001100;
		correct = 32'b00110011010011011001101000010101;
		#400 //2.7786455e+27 * 5.8045147e+34 = 4.787042e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110011101101101100001110010101;
		b = 32'b00110010000101010001000101001100;
		correct = 32'b11000001000111001110111100100100;
		#400 //-8.5106116e-08 * 8.676874e-09 = -9.808384
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110001110110100100010111100100;
		b = 32'b01010111000011011010111111101111;
		correct = 32'b10011010010001010010111111111101;
		#400 //-6.3525807e-09 * 155786770000000.0 = -4.077741e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100110011001111000101000110100;
		b = 32'b10101100101100110110000010110010;
		correct = 32'b01111001001001010011100011000101;
		#400 //-2.7335401e+23 * -5.0982213e-12 = 5.3617525e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010101111101000000110101101111;
		b = 32'b00101011110101001000010110100111;
		correct = 32'b00101001100100101111110110001110;
		#400 //9.857201e-26 * 1.5100602e-12 = 6.527687e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111111010001111111011001011001;
		b = 32'b10001011111000111010001111100110;
		correct = 32'b11110010111000001101111110111000;
		#400 //0.7811027 * -8.7683826e-32 = -8.908173e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011001001110100010011100000011;
		b = 32'b01000100111111000000010011110100;
		correct = 32'b01010011101111010001011110111001;
		#400 //3274827500000000.0 * 2016.1548 = 1624293600000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100110110011111000110001010100;
		b = 32'b10001111110000111101011110111101;
		correct = 32'b01010110100001111010011010000111;
		#400 //-1.4401546e-15 * -1.9311584e-29 = 74574650000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100110111100001000010110101101;
		b = 32'b11000101001010010100001100001001;
		correct = 32'b01100001001101011110001110001001;
		#400 //-5.6791692e+23 * -2708.1897 = 2.0970352e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010101011000011100111000001010;
		b = 32'b11110111111101101000000011010001;
		correct = 32'b10011100111010101000000100010101;
		#400 //15517190000000.0 * -9.999357e+33 = -1.5518188e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011110111000000001001110110000;
		b = 32'b00000101101011010000010111101110;
		correct = 32'b01011000101001011100010011010001;
		#400 //2.3725065e-20 * 1.627102e-35 = 1458117900000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100011110111010111111100100111;
		b = 32'b00000000100111010110110011011111;
		correct = 32'b01100010101101000001100001101111;
		#400 //2.4014719e-17 * 1.4457228e-38 = 1.6610873e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001001001110110111110100101011;
		b = 32'b11101010011000011101011010111111;
		correct = 32'b00011110010101001000011101000101;
		#400 //-767954.7 * -6.8255605e+25 = 1.125116e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111000000011011000010010000;
		b = 32'b10111001011110000001111000111011;
		correct = 32'b11001101000001011100111100111101;
		#400 //33200.562 * -0.00023662385 = -140309460.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101101111010100000001110011001;
		b = 32'b01001100001101111111101010111011;
		correct = 32'b01100001001000101100111110000011;
		#400 //9.05298e+27 * 48229100.0 = 1.8770783e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101101110001111111100111110100;
		b = 32'b00100100011110001100010111110000;
		correct = 32'b01001000110011011100100100100000;
		#400 //2.2734682e-11 * 5.3944087e-17 = 421449.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100011111110000010000001001101;
		b = 32'b11100010111100010111111111110110;
		correct = 32'b11000000100000111000001100011001;
		#400 //9.15424e+21 * -2.227443e+21 = -4.109753
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011011111111111001011001011100;
		b = 32'b00101001101110111001111100010101;
		correct = 32'b01110001101011100101111000111000;
		#400 //1.4388288e+17 * 8.3320646e-14 = 1.7268574e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001100110011110111011110010110;
		b = 32'b11010001001100001111010000101000;
		correct = 32'b00111011000101100001001001101100;
		#400 //-108772530.0 * -47500657000.0 = 0.0022899164
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011010111010100000010111101011;
		b = 32'b11110101111101101100111011000010;
		correct = 32'b10100100011100101011110101000011;
		#400 //3.2935826e+16 * -6.2573173e+32 = -5.2635696e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100110110000101000110001100100;
		b = 32'b10100110011011111111001100111010;
		correct = 32'b00111111110011111000111110111011;
		#400 //-1.3499507e-15 * -8.3249416e-16 = 1.6215738
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100100011101001011100111110111;
		b = 32'b11011111010101100111000001011100;
		correct = 32'b00000100100100100001010000101110;
		#400 //-5.3066584e-17 * -1.5451951e+19 = 3.4342967e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011101111100010011001000101110;
		b = 32'b11100101111110101100011110010000;
		correct = 32'b00110111011101100011011110001100;
		#400 //-2.1725006e+18 * -1.4803411e+23 = 1.4675676e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011101010011100011111100100010;
		b = 32'b01011110001101001100101010100001;
		correct = 32'b10111110100100100000010110101100;
		#400 //-9.288522e+17 * 3.2568505e+18 = -0.28519952
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001000001111111011000011011011;
		b = 32'b00111111101111101100101010001011;
		correct = 32'b00001000000000001001101010000100;
		#400 //5.7684864e-34 * 1.4905561 = 3.870023e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110111011001000101001111101001;
		b = 32'b01001010110100001011011001110101;
		correct = 32'b11101100000011000000011110010011;
		#400 //-4.6310374e+33 * 6839098.5 = -6.771415e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101001110000011101010101011101;
		b = 32'b00101011000101110011010101101001;
		correct = 32'b11111110001001000001010100011011;
		#400 //-2.9291283e+25 * 5.37201e-13 = -5.4525744e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111100110110111111100000100000;
		b = 32'b11011010010010100111110111000011;
		correct = 32'b01100010000010110000110001011101;
		#400 //-9.1371647e+36 * -1.4249055e+16 = 6.412471e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001101001110011001010001011001;
		b = 32'b00010101010011111011101100101111;
		correct = 32'b11110111011001001011001101111010;
		#400 //-194594190.0 * 4.195098e-26 = -4.638609e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101111100111100011100100110110;
		b = 32'b01011011001010111100010100101101;
		correct = 32'b11010011111010111100111101111001;
		#400 //-9.793559e+28 * 4.834902e+16 = -2025596300000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100100111000010010001000000101;
		b = 32'b10110011011110100001001011101100;
		correct = 32'b10110000111001100111011111001011;
		#400 //9.763583e-17 * -5.822487e-08 = -1.676875e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110101110110110101111111000011;
		b = 32'b01000000100000111001101100101101;
		correct = 32'b01110100110101010101110011101100;
		#400 //5.5617934e+32 * 4.1126924 = 1.3523485e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011111001010100001001011010010;
		b = 32'b10100010111001101011101001010111;
		correct = 32'b00111011101111001011001110111000;
		#400 //-3.6014468e-20 * -6.253892e-18 = 0.005758729
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110010110100100110100100000101;
		b = 32'b01100000110101000100010000010100;
		correct = 32'b01010001011111011100001100010000;
		#400 //8.335208e+30 * 1.2236298e+20 = 68118710000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011000111000011010010000111100;
		b = 32'b11001101100101111111101011000100;
		correct = 32'b10001010101111100000101000011100;
		#400 //5.832697e-24 * -318724220.0 = -1.8300137e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010101110000001110110110001111;
		b = 32'b01100101110000110100011000010110;
		correct = 32'b00101111011111001110110010111000;
		#400 //26515817000000.0 * 1.1526929e+23 = 2.3003366e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010001111111111101111001101111;
		b = 32'b01101011001010001111100101110111;
		correct = 32'b10100110010000011101001011001110;
		#400 //-137368560000.0 * 2.042776e+26 = -6.724602e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011010100101001010001010010001;
		b = 32'b11100101111100110010011111001001;
		correct = 32'b00110100000111000111110010010011;
		#400 //-2.091852e+16 * -1.4353362e+23 = 1.4573952e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100001100000110111111111111001;
		b = 32'b10100000101000110100001111100010;
		correct = 32'b01000000010011100011000100100111;
		#400 //-8.910779e-19 * -2.7658195e-19 = 3.22175
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010010111100010110001001010101;
		b = 32'b00101000000000101110000011100101;
		correct = 32'b00101010011011000001001101000000;
		#400 //1.5233479e-27 * 7.265216e-15 = 2.096769e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110100110000100011101001010010;
		b = 32'b00001000100000110011101110111110;
		correct = 32'b11101011101111010111000100111111;
		#400 //-3.617775e-07 * 7.898321e-34 = -4.5804354e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111000010010011011011010011010;
		b = 32'b01111011110000011100110001011111;
		correct = 32'b00111100000001010011101001001001;
		#400 //1.6364926e+34 * 2.0125169e+36 = 0.008131572
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000001001101011001100011100000;
		b = 32'b00010110111000111110110011000101;
		correct = 32'b01101001110010111111011100111101;
		#400 //11.349823 * 3.682325e-25 = 3.0822436e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101011011001110001101001001111;
		b = 32'b01000110010101001101100100011110;
		correct = 32'b11100100100010101111101001001111;
		#400 //-2.793861e+26 * 13622.279 = -2.0509499e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101010011110101010000100101111;
		b = 32'b01001111100011011011000101011001;
		correct = 32'b10011010011000100110100011010111;
		#400 //-2.2260382e-13 * 4754420000.0 = -4.6820394e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111100101110011011101111110110;
		b = 32'b01111010110101111001000111110001;
		correct = 32'b10000001010111001001000110000110;
		#400 //-0.022672635 * 5.5965193e+35 = -4.0512026e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100110001101000010000011011101;
		b = 32'b10110011000111101001101100000011;
		correct = 32'b11110010100100010101111010100011;
		#400 //2.1265805e+23 * -3.6928224e-08 = -5.758686e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100110100111011000011101001010;
		b = 32'b01111101100110100100000110011011;
		correct = 32'b00101000100000101011011100011010;
		#400 //3.719536e+23 * 2.563022e+37 = 1.4512307e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111000111010001100110000111001;
		b = 32'b00100111100111011101110101110101;
		correct = 32'b11010000101111001100000111000000;
		#400 //-0.000111006615 * 4.381636e-15 = -25334514000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101011111101110000100001100000;
		b = 32'b01001101001000001101010100110101;
		correct = 32'b10011110010001001001101001010001;
		#400 //-1.755273e-12 * 168645460.0 = -1.04080655e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001011011111000001000010010111;
		b = 32'b01001110110001001110101000000010;
		correct = 32'b00111100001000111101100101111111;
		#400 //16519319.0 * 1651835100.0 = 0.010000586
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010011110110101011111000111100;
		b = 32'b00100001010001000001001100010111;
		correct = 32'b00110010000011101100110001011110;
		#400 //5.5218522e-27 * 6.643265e-19 = 8.311956e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111100111100000100110110001110;
		b = 32'b01111100001100100011000000111000;
		correct = 32'b11000000001011001001111010010101;
		#400 //-9.981794e+36 * 3.7008273e+36 = -2.697179
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111010001010010100011001100010;
		b = 32'b10101001001011110010101110111010;
		correct = 32'b11010000011101110110001000110011;
		#400 //0.0006457326 * -3.8895733e-14 = -16601632000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010101101010101001011001000000;
		b = 32'b11010001110010101111100111000001;
		correct = 32'b11000011010101110010011001110110;
		#400 //23445287000000.0 * -108971700000.0 = -215.15024
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101000001101100011110110010101;
		b = 32'b01000011100010111101100010110011;
		correct = 32'b00100100001001101100110110000111;
		#400 //1.0116383e-14 * 279.69296 = 3.61696e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000101011000111010000101110000;
		b = 32'b11001101100011101011110000001110;
		correct = 32'b00110111010011000010000111010101;
		#400 //-3642.0898 * -299336130.0 = 1.2167225e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011001011111111010010101101111;
		b = 32'b00011101000001001100111010010010;
		correct = 32'b00111011111101100110010010100111;
		#400 //1.32166e-23 * 1.7576849e-21 = 0.007519323
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000111011111110111101100101100;
		b = 32'b10110111000011111101101011011110;
		correct = 32'b10001111111000110101001011000110;
		#400 //1.9220265e-34 * -8.574423e-06 = -2.2415811e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101001111001001100111110011000;
		b = 32'b10010110011001111000101011100010;
		correct = 32'b11010010111111001111101011011001;
		#400 //1.0161246e-13 * -1.8703855e-25 = -543270140000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011111000100001011110101010011;
		b = 32'b10000001110111101011101110000000;
		correct = 32'b01011100101001100101101110100111;
		#400 //-3.064979e-20 * -8.181897e-38 = 3.7460495e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100110111001111000000000010000;
		b = 32'b00101101101000001100010010000001;
		correct = 32'b00111000101110000101000011100010;
		#400 //1.6063556e-15 * 1.827716e-11 = 8.788869e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101010100100011110010010110000;
		b = 32'b01101110110001101100011011111000;
		correct = 32'b10111011001110111110010001100111;
		#400 //-8.8187095e+25 * 3.0759285e+28 = -0.0028670074
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010110000100100011000000101101;
		b = 32'b10000111011111011000011111110111;
		correct = 32'b11001110000100111001110010011101;
		#400 //1.1808988e-25 * -1.9073561e-34 = -619128640.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111101001100011100100101110011;
		b = 32'b01001101010010000110001011100111;
		correct = 32'b01101111011000110010000011100110;
		#400 //1.4769959e+37 * 210120300.0 = 7.029287e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110010110101010010100110000100;
		b = 32'b01001001110101001001110000011011;
		correct = 32'b00101000100000000101010100100011;
		#400 //2.4815343e-08 * 1741699.4 = 1.4247777e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101111101100011101011101000101;
		b = 32'b00010010110011100000110110011100;
		correct = 32'b01011100010111001111001011111011;
		#400 //3.234907e-10 * 1.3003783e-27 = 2.4876662e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000000110101001001011001000011;
		b = 32'b11110111010101000001011111110100;
		correct = 32'b00001001000000000100110000111010;
		#400 //-6.6433425 * -4.3017686e+33 = 1.5443281e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111110011111110100000110101;
		b = 32'b11010100100001110000110111101011;
		correct = 32'b00100010110001010000110000011110;
		#400 //-2.4784453e-05 * -4640432700000.0 = 5.3409787e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101110110001100101101010101011;
		b = 32'b10110101100111110001100111011010;
		correct = 32'b10111000100111111001010001111011;
		#400 //9.0201034e-11 * -1.1853947e-06 = -7.6093675e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111110111110011101100110111110;
		b = 32'b01110111001101101001101010110010;
		correct = 32'b11000111001011110010001100111000;
		#400 //-1.6605418e+38 * 3.7036548e+33 = -44835.22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101010010001011110010110101010;
		b = 32'b11010001000101100100111110000111;
		correct = 32'b00011000101010001000010111110000;
		#400 //-1.7576796e-13 * -40348710000.0 = 4.3562224e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011110000101111010010111111110;
		b = 32'b01100001001010100110111111100000;
		correct = 32'b00111100011000111100011101110100;
		#400 //2.7318548e+18 * 1.965005e+20 = 0.013902534
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100001100100100001100011011001;
		b = 32'b10111010001011111110001000101000;
		correct = 32'b01100110110101001010010101001010;
		#400 //-3.368769e+20 * -0.000670942 = 5.0209537e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010100011011011011011100011010;
		b = 32'b00111010011100100011010110111111;
		correct = 32'b10011001011110110011111111011000;
		#400 //-1.2001553e-26 * 0.0009239576 = -1.2989289e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110101110010101110111001111111;
		b = 32'b00100101111111001001101111110000;
		correct = 32'b11001111010011011010011111011001;
		#400 //-1.5119584e-06 * 4.38207e-16 = -3450329300.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001001010110110010101011010011;
		b = 32'b11011010001000100101111010100011;
		correct = 32'b10101110101011001100011001100011;
		#400 //897709.2 * -1.142575e+16 = -7.856895e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111101011011101111001000000011;
		b = 32'b11101100011110010010001101101000;
		correct = 32'b10010000011101011000011010111101;
		#400 //0.05833627 * -1.2047589e+27 = -4.842153e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111011101110001101000100000011;
		b = 32'b01111111110110001000111001110100;
		correct = 32'b01111111110110001000111001110100;
		#400 //0.0056401505 * nan = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100001111000111010110001101101;
		b = 32'b01010011000000011111111011000111;
		correct = 32'b01001110011000000010110111011010;
		#400 //5.2497944e+20 * 558325240000.0 = 940275300.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101101110110110101100010001100;
		b = 32'b11100100010110101011001111101100;
		correct = 32'b11001001000000000110000001011010;
		#400 //8.485533e+27 * -1.613742e+22 = -525829.6
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010010110111010001010110000111;
		b = 32'b01111101111000001110001010111101;
		correct = 32'b00010100011110111010110000100100;
		#400 //474774470000.0 * 3.7365545e+37 = 1.270621e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110010001110101110001100000;
		b = 32'b11101100000111101010010111110011;
		correct = 32'b10010001101000001101100011111100;
		#400 //0.19468832 * -7.671758e+26 = -2.5377276e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011100101101101011000111011010;
		b = 32'b00110111111110000111010010110101;
		correct = 32'b10100100001111000011110111111001;
		#400 //-1.2089723e-21 * 2.961825e-05 = -4.0818495e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000011001101000111110000111001;
		b = 32'b00001010110101011100111010111001;
		correct = 32'b01110111110110000001101000011010;
		#400 //180.48524 * 2.0588914e-32 = 8.766137e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000000001110100110000001100011;
		b = 32'b10011011001001101010010001001011;
		correct = 32'b01100100100011110010100010010110;
		#400 //-2.912133 * -1.3784284e-22 = 2.1126471e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100111000111011111110000001100;
		b = 32'b10111010010110101111101111110001;
		correct = 32'b11101100001110001011000001111011;
		#400 //7.46061e+23 * -0.0008353582 = -8.93103e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010101001101110101100110101100;
		b = 32'b11110011101100011011011100000010;
		correct = 32'b10100001000001000000111100010110;
		#400 //12599735000000.0 * -2.8160046e+31 = -4.4743306e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111001001100101100101110111111;
		b = 32'b00111111010101100010010001100011;
		correct = 32'b11111001010101011011111010100101;
		#400 //-5.802258e+34 * 0.8364927 = -6.9364123e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001001010101001111101011010110;
		b = 32'b01011110010101011100000110010000;
		correct = 32'b10101010011111110001001000000000;
		#400 //-872365.4 * 3.8506876e+18 = -2.2654795e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010110011111111001100000101011;
		b = 32'b10111100001010001100011101001111;
		correct = 32'b01011001110000011101011100011110;
		#400 //-70257255000000.0 * -0.010301425 = 6820149300000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001010111000111100101010110011;
		b = 32'b11010101010101100111110110011011;
		correct = 32'b00110101000001111111000000001000;
		#400 //-7464281.5 * -14739685000000.0 = 5.064071e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101000101010011100111010100100;
		b = 32'b10011100011000101010001001101001;
		correct = 32'b11001011101111111100111100111101;
		#400 //1.8852385e-14 * -7.498704e-22 = -25140858.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000110110110010100101111001010;
		b = 32'b11100110000110101110001011010001;
		correct = 32'b10100000001100111001001110011001;
		#400 //27813.895 * -1.8285712e+23 = -1.5210726e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000011000111001010111100111100;
		b = 32'b00110011010111010000001110101011;
		correct = 32'b01001111001101010111110010101110;
		#400 //156.68451 * 5.145891e-08 = 3044847000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000101101000001100000101111000;
		b = 32'b10100000000111100001011101111100;
		correct = 32'b00100101000000100010100000101100;
		#400 //-1.5117397e-35 * -1.3390891e-19 = 1.1289313e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101000001101111101111100011001;
		b = 32'b10111101100111010000011010011000;
		correct = 32'b00101010000101011110001000100100;
		#400 //-1.0206917e-14 * -0.07667273 = 1.3312317e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011100101010100111011101010110;
		b = 32'b11100101100110010010001110111000;
		correct = 32'b10110110100011100111101101110110;
		#400 //3.8385566e+17 * -9.039762e+22 = -4.2463025e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110001110110011110111110011110;
		b = 32'b10001100000011000101001010100000;
		correct = 32'b01100101010001101100110000100111;
		#400 //-6.3427725e-09 * -1.0810072e-31 = 5.8674657e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100011101110000011010011101011;
		b = 32'b11010101001000010010001100011011;
		correct = 32'b10001110000100100101001101001111;
		#400 //1.9971732e-17 * -11073259000000.0 = -1.8036001e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110100101111001001101010100111;
		b = 32'b11011110101100010000001110100111;
		correct = 32'b11010101100010000110000101110100;
		#400 //1.1954206e+32 * -6.377611e+18 = -18744017000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100100011011110111111110110011;
		b = 32'b00001000111110101111101000000010;
		correct = 32'b11011010111101000100101011100001;
		#400 //-5.193303e-17 * 1.5105104e-33 = -3.4381112e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110010100110111100000100110011;
		b = 32'b01111000100100011001000111100100;
		correct = 32'b00111001100010001111010010011101;
		#400 //6.170079e+30 * 2.3620064e+34 = 0.00026122193
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111111010101110000001101011011;
		b = 32'b11001000000110010100111100100001;
		correct = 32'b11110110101100111000010010000000;
		#400 //2.8580144e+38 * -156988.52 = -1.8205245e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000011011001101011111010011100;
		b = 32'b00111101011110011001111001000100;
		correct = 32'b11000101011011001010010011010001;
		#400 //-230.74457 * 0.06094195 = -3786.301
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000111000001111101000101100010;
		b = 32'b11011100011001101111111011101010;
		correct = 32'b00101010000101101000010100000011;
		#400 //-34769.383 * -2.600781e+17 = 1.3368824e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010100001011110111110011001000;
		b = 32'b11000011100011000001111110110101;
		correct = 32'b11010000001000000100110111001000;
		#400 //3014851000000.0 * -280.2477 = -10757808000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111001000010100100100111101101;
		b = 32'b10111100010111110011111010111011;
		correct = 32'b11111100000111101001010000101011;
		#400 //4.487727e+34 * -0.013625796 = -3.2935524e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110110101110001010111011011001;
		b = 32'b01110100100000100000100110010001;
		correct = 32'b00000001101101011100101000011010;
		#400 //5.5039823e-06 * 8.242097e+31 = 6.67789e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001110111111000100111110100101;
		b = 32'b10010011100010000110011110111111;
		correct = 32'b10111010111011001100001110000110;
		#400 //6.219949e-30 * -3.443353e-27 = -0.0018063642
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010111011100000001011110100101;
		b = 32'b11000110111011001100101000101101;
		correct = 32'b00010000000000011100100100001000;
		#400 //-7.7578026e-25 * -30309.088 = 2.5595633e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010101011110011111001010010010;
		b = 32'b01010110110001100101111000101110;
		correct = 32'b10111110001000010100100001010111;
		#400 //-17176264000000.0 * 109053900000000.0 = -0.15750252
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100110011000111001111111010110;
		b = 32'b01100000111101001011110100010110;
		correct = 32'b10000100111011100001100100100111;
		#400 //-7.8973064e-16 * 1.4108221e+20 = -5.597663e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110100010100000000010110001100;
		b = 32'b01000101101000100111001000110011;
		correct = 32'b10101110001000111110100101010100;
		#400 //-1.9373527e-07 * 5198.275 = -3.7269146e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011101001110000110101101111010;
		b = 32'b01000110000101010010110010111000;
		correct = 32'b11010110100111100011111000000100;
		#400 //-8.305531e+17 * 9547.18 = -86994600000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010010101101111111111000011000;
		b = 32'b00111101110000110111100011110101;
		correct = 32'b10010100011100001111011100100000;
		#400 //-1.1611563e-27 * 0.09544555 = -1.216564e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111101110000100010110011010101;
		b = 32'b11100001101100001111000011010001;
		correct = 32'b01011011100011000111011110101110;
		#400 //-3.2262877e+37 * -4.0799745e+20 = 7.907617e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000111101000011010111100101;
		b = 32'b00010100011000100110111000011010;
		correct = 32'b11011100000010100000110100011100;
		#400 //-1.7768654e-09 * 1.1431798e-26 = -1.5543184e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000001111001011101011100000011;
		b = 32'b00011101110100000100011011000000;
		correct = 32'b10100011100011010100000010010100;
		#400 //-8.442984e-38 * 5.5130295e-21 = -1.53146e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101011001110111010001000011000;
		b = 32'b10101100001111011111010001101011;
		correct = 32'b00111110011111001101111100001001;
		#400 //-6.6660696e-13 * -2.6994195e-12 = 0.24694456
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011100001101110111111101101110;
		b = 32'b00100011001101100011000011000101;
		correct = 32'b00111000100000001110101100011111;
		#400 //6.071432e-22 * 9.876567e-18 = 6.14731e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110010111000010111010010111001;
		b = 32'b01101110100111101000100101011010;
		correct = 32'b01000011101101100000011110011100;
		#400 //8.93123e+30 * 2.453234e+28 = 364.05945
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000101100100001111011110000100;
		b = 32'b00101100000110001010001011011111;
		correct = 32'b11011000111100110010001100010100;
		#400 //-4638.9395 * 2.169091e-12 = -2138655900000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011000110101011011010000001101;
		b = 32'b01010000010001010110101001101111;
		correct = 32'b01001000000010101000111101111101;
		#400 //1879754300000000.0 * 13248347000.0 = 141885.95
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110000111111111111010110011000;
		b = 32'b10110111111000100010000100010010;
		correct = 32'b10111000100100001110001010100100;
		#400 //1.8623494e-09 * -2.6956699e-05 = -6.90867e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101110001111001001000011110010;
		b = 32'b11110100110100100011010010010111;
		correct = 32'b10111000111001011010010110000010;
		#400 //1.4589602e+28 * -1.3323352e+32 = -0.00010950399
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001010100011001001010111110101;
		b = 32'b00001110011000111100101110010011;
		correct = 32'b00111011100111011111111000011011;
		#400 //1.3537917e-32 * 2.8077928e-30 = 0.0048215515
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010101010010101111011000011001;
		b = 32'b01001001011110000110101011000010;
		correct = 32'b01001011010100010010100000100001;
		#400 //13947396000000.0 * 1017516.1 = 13707297.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010011111100001101111011110000;
		b = 32'b01000111011011010101011010001000;
		correct = 32'b11001100000000011110011111000011;
		#400 //-2069064800000.0 * 60758.53 = -34053900.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001001010001110000010101101111;
		b = 32'b00001100000000111010100100110111;
		correct = 32'b00111100110000010111110010111001;
		#400 //2.3956309e-33 * 1.0142794e-31 = 0.023619043
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011111111000111101010100001011;
		b = 32'b00010101000100100000100011101110;
		correct = 32'b11001010010001111011001000010010;
		#400 //-9.649069e-20 * 2.949151e-26 = -3271812.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011110001000111000111100010001;
		b = 32'b00110110000001110100000001111000;
		correct = 32'b11100111100110101100101000001110;
		#400 //-2.9464144e+18 * 2.0154093e-06 = -1.4619434e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111101101100100110001000110011;
		b = 32'b00011101011000100100100111100101;
		correct = 32'b01011111110010011100111000011010;
		#400 //0.08710136 * 2.9949054e-21 = 2.9083178e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001011100100101010100011110000;
		b = 32'b00011011011000010010101011110011;
		correct = 32'b10101111101001101011110111111000;
		#400 //-5.6491343e-32 * 1.8625441e-22 = -3.0330205e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111000001010011011110001101011;
		b = 32'b11011100010000111111011010011001;
		correct = 32'b01011011010111011011110011010001;
		#400 //-1.3770621e+34 * -2.2063503e+17 = 6.2413576e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011011000101111001010111111001;
		b = 32'b10100010101101110001001011011110;
		correct = 32'b01110111110100111111100000011001;
		#400 //-4.266762e+16 * -4.9622226e-18 = 8.5984895e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001010011000110000011011011001;
		b = 32'b10001101010011100101110000001100;
		correct = 32'b11111100100011001101000111000011;
		#400 //3719606.2 * -6.358945e-31 = -5.849408e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100001101000100010110111100001;
		b = 32'b10000011101010110110010111101110;
		correct = 32'b01011101011100100011101100001000;
		#400 //-1.0989691e-18 * -1.0073879e-36 = 1.0909096e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110101000111110011110101100111;
		b = 32'b10111101001101011100000000111011;
		correct = 32'b01110111011000000100101011101111;
		#400 //-2.018605e+32 * -0.04437278 = 4.5491966e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011111011010101000000101010110;
		b = 32'b10100100110011110111010001001111;
		correct = 32'b01111010000100001011000011000100;
		#400 //-1.6897882e+19 * -8.9968974e-17 = 1.87819e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110010100111110110001100101001;
		b = 32'b10111010101101000010110100011100;
		correct = 32'b10110111011000100111011001101000;
		#400 //1.8555129e-08 * -0.0013746354 = -1.3498218e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100101110011111011011011111011;
		b = 32'b10101000110110010110101110010000;
		correct = 32'b11111100011101001001001010001011;
		#400 //1.2261316e+23 * -2.4138487e-14 = -5.0795707e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000011101001001000001100000000;
		b = 32'b01100101000100111101110010001110;
		correct = 32'b10011110000011100110100111100100;
		#400 //-329.02344 * 4.3641024e+22 = -7.539315e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111111000000101001100110010000;
		b = 32'b11000000000000101011101010001101;
		correct = 32'b10111110011111111011111101100111;
		#400 //0.5101557 * -2.0426362 = -0.24975358
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111011111111000001101000110010;
		b = 32'b10110111100010010110000101111011;
		correct = 32'b11000011111010101110001101010100;
		#400 //0.0076935524 * -1.6377066e-05 = -469.776
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100010101011100111100001111011;
		b = 32'b10001000010100101000011000101011;
		correct = 32'b11011001110101000010100010010101;
		#400 //4.729036e-18 * -6.335229e-34 = -7464664400000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101100100011100001010101001110;
		b = 32'b01101010111001111000111101010000;
		correct = 32'b01000001000111010001010001011011;
		#400 //1.3741446e+27 * 1.3996932e+26 = 9.81747
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110000100100011001100101110;
		b = 32'b10010000101101110110000001101110;
		correct = 32'b01100100110011000001100110011001;
		#400 //-2.1785486e-06 * -7.2329346e-29 = 3.0119842e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110101101001011110100111101110;
		b = 32'b01101110001110001110101000011000;
		correct = 32'b01000110111001011011000111101111;
		#400 //4.2064143e+32 * 1.4307061e+28 = 29400.967
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001001011111101101000110101110;
		b = 32'b00011011100100010000100000010001;
		correct = 32'b01101101011000001110010100010101;
		#400 //1043738.9 * 2.399345e-22 = 4.350099e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100001101101000001111000001111;
		b = 32'b00101011011100010111011110101001;
		correct = 32'b11110101101111101111010100101010;
		#400 //-4.153225e+20 * 8.578646e-13 = -4.841352e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111001110000110000011100101011;
		b = 32'b01000110010110001001000110111001;
		correct = 32'b10110010111001101000100101101001;
		#400 //-0.0003719864 * 13860.431 = -2.6838011e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010100100100000001101111100011;
		b = 32'b01111000000001100100011111011011;
		correct = 32'b00011100000010010101111001011001;
		#400 //4951545000000.0 * 1.0894143e+34 = 4.545144e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110100110100000001001001010000;
		b = 32'b11100011101111001100100100011111;
		correct = 32'b11010000100011010001001110000001;
		#400 //1.31881e+32 * -6.9649604e+21 = -18934925000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110000111111111100110000101010;
		b = 32'b11111110100001110010001111101110;
		correct = 32'b10110001111100100100100000110101;
		#400 //6.3332397e+29 * -8.981617e+37 = -7.051336e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111011101100100100000101110101;
		b = 32'b11001100110001000100010111010111;
		correct = 32'b11101110011010001000000000001001;
		#400 //1.851113e+36 * -102903480.0 = -1.7988827e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001111001010100110101000110001;
		b = 32'b01011101010101000101011100111101;
		correct = 32'b10110001010011010111010000100100;
		#400 //-2859086000.0 * 9.562978e+17 = -2.9897445e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111011100100101101001000110011;
		b = 32'b11000000100001000000000000100011;
		correct = 32'b01111010100011100101111100010011;
		#400 //-1.5246774e+36 * -4.1250167 = 3.6961724e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010011111110110110110010111111;
		b = 32'b10000011111110110001110101001111;
		correct = 32'b01001111100000000010100001111110;
		#400 //-6.346854e-27 * -1.4759183e-36 = 4300274700.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110111101101111010101111111011;
		b = 32'b10111001001111111100111111000110;
		correct = 32'b10111101111101010010001011100001;
		#400 //2.1895385e-05 * -0.00018292581 = -0.11969543
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101010100010001111010011101000;
		b = 32'b11001100100101000101010001100110;
		correct = 32'b10011101011011000101111100011001;
		#400 //2.432839e-13 * -77767470.0 = -3.1283504e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000010010110001101000100110111;
		b = 32'b00000110010110000011110101011110;
		correct = 32'b10111011100000000101011110000100;
		#400 //-1.5929215e-37 * 4.067017e-35 = -0.0039166827
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111001101110111100000001010011;
		b = 32'b11000011111000101000101000111111;
		correct = 32'b00110101010101000010101011000011;
		#400 //-0.00035810712 * -453.08005 = 7.903838e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101111101010100011001010100111;
		b = 32'b01001000011011010110110110000110;
		correct = 32'b10100110101101111000001011011010;
		#400 //-3.095881e-10 * 243126.1 = -1.2733643e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001100110001110010101101100011;
		b = 32'b10110001000001100000000000010110;
		correct = 32'b00011011001111100100000000111111;
		#400 //-3.0686917e-31 * -1.9499615e-09 = 1.5737191e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011010111110011110100011010000;
		b = 32'b11100101111100010101010110000100;
		correct = 32'b10110100100001001000110001011010;
		#400 //3.5171625e+16 * -1.4245848e+23 = -2.4689035e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101110100010001111000000010101;
		b = 32'b10111011001011101100011111101001;
		correct = 32'b01110010110010001001001001010011;
		#400 //-2.1190101e+28 * -0.0026669449 = 7.945459e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001010110110001000010111110000;
		b = 32'b00100010100110100101000101001011;
		correct = 32'b11100111101100111001100011010101;
		#400 //-7095032.0 * 4.1827856e-18 = -1.6962457e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000111000101101011010110000100;
		b = 32'b10100100000111111000000101101100;
		correct = 32'b10100010011100011110000111001000;
		#400 //1.1338088e-34 * -3.4587254e-17 = -3.2781118e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100000111001111100110011101100;
		b = 32'b10111100010000000101010010111110;
		correct = 32'b10100100000110100100010010000111;
		#400 //3.9268528e-19 * -0.011738954 = -3.3451472e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110101001101010101111001000010;
		b = 32'b01001101011111011010111011011000;
		correct = 32'b01100111001101110000011001010100;
		#400 //2.299115e+32 * 266005890.0 = 8.643098e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110110001110001001110010110100;
		b = 32'b01111001111111001100111010001001;
		correct = 32'b00111011101110101111000110101000;
		#400 //9.360947e+32 * 1.6408098e+35 = 0.005705077
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001110111010101101000110101011;
		b = 32'b01011000101110111101111101111100;
		correct = 32'b10110101100111111111110000100000;
		#400 //-1969804700.0 * 1652548300000000.0 = -1.1919801e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110100010111111110001011101;
		b = 32'b11011011100110100010000000100011;
		correct = 32'b10100010011010001000001110011110;
		#400 //0.27340975 * -8.676496e+16 = -3.151154e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111000111100010011010000110010;
		b = 32'b11000101001100011111001111111000;
		correct = 32'b10110011001011010111111011101100;
		#400 //0.00011501498 * -2847.248 = -4.0395136e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001101000000100010100000000101;
		b = 32'b00110011011110101000100001110101;
		correct = 32'b01011001000001001111111100011011;
		#400 //136478800.0 * 5.8331768e-08 = 2339699300000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101010100111010110111111001001;
		b = 32'b11110101100010101111101000000100;
		correct = 32'b10110100100100010000000010000101;
		#400 //9.516462e+25 * -3.523476e+32 = -2.7008733e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010001110111110000001001000100;
		b = 32'b00100011111111001101100001010011;
		correct = 32'b11101101011000011100101010100010;
		#400 //-119726965000.0 * 2.7413512e-17 = -4.3674435e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000110101110111011010110001111;
		b = 32'b10000000001111101111011011000000;
		correct = 32'b01000110001111101100110001010100;
		#400 //-7.060836e-35 * -5.782318e-39 = 12211.082
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000101000011001100100110001011;
		b = 32'b10000101001011000001110100101000;
		correct = 32'b10111111010100010110011110111011;
		#400 //6.619786e-36 * -8.092756e-36 = -0.81798905
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010111010011110111010111111110;
		b = 32'b11011001100100000101110111001000;
		correct = 32'b00111101001101111111000100010111;
		#400 //-228105680000000.0 * -5079439000000000.0 = 0.044907656
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111001011110111100001111110100;
		b = 32'b11000000011101001011110111100111;
		correct = 32'b00111000100000111010110001100001;
		#400 //-0.00024010224 * -3.8240907 = 6.278675e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001010111100111000000000000001;
		b = 32'b10101110001010010000011010001000;
		correct = 32'b11011100001110000110010111110001;
		#400 //7979008.5 * -3.8431952e-11 = -2.0761393e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101110011011111111010011110011;
		b = 32'b11110100100101100001010001000010;
		correct = 32'b00111001010011001010011110111011;
		#400 //-1.8565761e+28 * -9.512395e+31 = 0.0001951744
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100000000110011011110000001000;
		b = 32'b10011100111001100000100010111110;
		correct = 32'b01000010101010110001011001111001;
		#400 //-1.3021818e-19 * -1.5222383e-21 = 85.54389
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000100001001011010100101100010;
		b = 32'b10000100001111111001010111111101;
		correct = 32'b10111111010111010101110000010001;
		#400 //1.9473434e-36 * -2.2520813e-36 = -0.8646861
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100100001111010101111101010101;
		b = 32'b01011100001011011111100110000000;
		correct = 32'b01000111100010110101010000101001;
		#400 //1.3973216e+22 * 1.95878e+17 = 71336.32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011001110111101110010011010101;
		b = 32'b00100101001111110011100100011101;
		correct = 32'b00110100000101010011001100011011;
		#400 //2.3046687e-23 * 1.658596e-16 = 1.3895298e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001110111111111001100100110111;
		b = 32'b01001000100000110111110010010101;
		correct = 32'b00000101111110001101001000011101;
		#400 //6.3009894e-30 * 269284.66 = 2.3398991e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110100010011011100111111100100;
		b = 32'b01000000101011000000101000111001;
		correct = 32'b11110011000110010010000001111110;
		#400 //-6.522445e+31 * 5.376248 = -1.2131965e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000100101110111101010101001010;
		b = 32'b00010101111111011001110100000001;
		correct = 32'b00101110001111011001100111001111;
		#400 //4.4159364e-36 * 1.02433595e-25 = 4.3110234e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001100001011000111100010110100;
		b = 32'b11111110100101010100110000101100;
		correct = 32'b10001101000100111101111000111111;
		#400 //45212370.0 * -9.922524e+37 = -4.556539e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010000101110110110100010110111;
		b = 32'b11101110001000010000111100101010;
		correct = 32'b10100010000101001111000011110011;
		#400 //25153616000.0 * -1.2461355e+28 = -2.0185298e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011010110010000001010111000110;
		b = 32'b00101010000111101110110101100011;
		correct = 32'b00110000001000010010011000000001;
		#400 //8.275324e-23 * 1.4115579e-13 = 5.8625466e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100000001010101100010100001110;
		b = 32'b11110101101011001010000000000010;
		correct = 32'b10101001111111010011111110100111;
		#400 //4.9221028e+19 * -4.3765645e+32 = -1.1246499e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000111101000001100010000101000;
		b = 32'b01100101101111110101011110011010;
		correct = 32'b10100001010101110001011110000111;
		#400 //-82312.31 * 1.12948495e+23 = -7.287597e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101001010001111011000110010111;
		b = 32'b01000111000001110100110000110100;
		correct = 32'b11100001101111001110110000110011;
		#400 //-1.508843e+25 * 34636.203 = -4.3562598e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011111001000101010010001001001;
		b = 32'b01010011011100011001110000001001;
		correct = 32'b11001011001011000101010000101110;
		#400 //-1.1719572e+19 * 1037704950000.0 = -11293742.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111001011001001001010011001;
		b = 32'b10111010101111111010111100101100;
		correct = 32'b11001011111001100111100111010011;
		#400 //44178.598 * -0.0014624349 = -30208934.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010000111101011100101101100011;
		b = 32'b01001011000101000101111001111110;
		correct = 32'b01000101010101000000110011010111;
		#400 //32989977000.0 * 9723518.0 = 3392.8025
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001101111111010100010001101011;
		b = 32'b00101010100110001000100100010101;
		correct = 32'b01100010110101001000011101101011;
		#400 //531139940.0 * 2.7095744e-13 = 1.9602338e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010011111001000110100010000111;
		b = 32'b00000001010111010000100001001010;
		correct = 32'b01010010000001000100010101111011;
		#400 //5.7658364e-27 * 4.0597236e-38 = 142025340000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110000101100010011110111101101;
		b = 32'b11001010000001111101100001010000;
		correct = 32'b01100110001001110000000110011011;
		#400 //-4.388297e+29 * -2225684.0 = 1.971662e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110101111100111101110111110111;
		b = 32'b11111011110110110001001101110101;
		correct = 32'b00111001100011100111110000010110;
		#400 //-6.1827643e+32 * -2.2750153e+36 = 0.00027176802
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111001011010110010011001000001;
		b = 32'b11000101100110111001111010111000;
		correct = 32'b10110011010000010110101000001101;
		#400 //0.00022425597 * -4979.84 = -4.5032767e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101001000001001000000010001111;
		b = 32'b01111000101011000010101101001110;
		correct = 32'b10101111110001010000010011001111;
		#400 //-1.0011582e+25 * 2.7936043e+34 = -3.5837508e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111111111100011011101100100101;
		b = 32'b11011101010100011110000001011100;
		correct = 32'b01111111111100011011101100100101;
		#400 //nan * -9.451993e+17 = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010011101011100011011000100110;
		b = 32'b00000010110101111010011111000011;
		correct = 32'b11010000010011101100110110001100;
		#400 //-4.397717e-27 * 3.1687701e-37 = -13878309000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111101110010101011001011000001;
		b = 32'b01011100000111111011001001001110;
		correct = 32'b00100001001000100111011101111111;
		#400 //0.09897376 * 1.7980228e+17 = 5.5045887e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101001111110111011001001100001;
		b = 32'b01011000110101010100001011100111;
		correct = 32'b00010000100101110001000110101110;
		#400 //1.1177583e-13 * 1875866600000000.0 = 5.958624e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011011011101010011000001011010;
		b = 32'b11010001101011100110101001001010;
		correct = 32'b00001001001100111111000010000001;
		#400 //-2.0281548e-22 * -93638440000.0 = 2.1659426e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010101111110100111010100110010;
		b = 32'b00101000100111011110001100110000;
		correct = 32'b10101100110010110000110000010010;
		#400 //-1.011591e-25 * 1.7529028e-14 = -5.770947e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010110000110001101011010011000;
		b = 32'b01110011011000101010010010111000;
		correct = 32'b10100010001011001010001010010001;
		#400 //-42011860000000.0 * 1.7956543e+31 = -2.3396409e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110001010011110100110000111100;
		b = 32'b11001000010011010110110010110011;
		correct = 32'b00101000100000010010101011001100;
		#400 //-3.0165799e-09 * -210354.8 = 1.4340437e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111010001000110110001110101;
		b = 32'b00110001101000000010110101011001;
		correct = 32'b01010101000111001111011100010100;
		#400 //50284.457 * 4.6617683e-09 = 10786563000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111001111111100010110011110;
		b = 32'b10100000101111000010111011100010;
		correct = 32'b11100110000000100111000011101010;
		#400 //49093.617 * -3.1879463e-19 = -1.5399763e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011100001100110100111101010010;
		b = 32'b00100011101101110100001010001001;
		correct = 32'b10110111111110100111101101101001;
		#400 //-5.932865e-22 * 1.9869078e-17 = -2.985979e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011110110011001111000110011;
		b = 32'b10110001011010110111111001000010;
		correct = 32'b01011001111011001001000101110101;
		#400 //-28523622.0 * -3.426877e-09 = 8323503300000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011110111011011001010100001000;
		b = 32'b01001001000010001111110011110100;
		correct = 32'b10010101010111011111111001101101;
		#400 //-2.5154989e-20 * 561103.25 = -4.48313e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010100111111011110011001011111;
		b = 32'b00100100110001001000110000011001;
		correct = 32'b11101111101001010101100110111010;
		#400 //-8723933700000.0 * 8.5238785e-17 = -1.02347e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011010110110111101011110101110;
		b = 32'b10111000111110110000011000111101;
		correct = 32'b01100001011000000011001100110111;
		#400 //-3.0940081e+16 * -0.00011969775 = 2.5848507e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101000101011001100000000000110;
		b = 32'b11010010100011111111111000001011;
		correct = 32'b01010101100110011001000001010100;
		#400 //-6.526314e+24 * -309221230000.0 = 21105645000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001101000110101011110110001100;
		b = 32'b00110000101000111100100000111111;
		correct = 32'b01011011111100011101111000000010;
		#400 //162257090.0 * 1.1916724e-09 = 1.3615914e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000100000010111101000101001110;
		b = 32'b00000110101111011000110110010010;
		correct = 32'b11111100101111001101010001111110;
		#400 //-559.2704 * 7.130192e-35 = -7.843693e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010100011011001101010010101010;
		b = 32'b00011111010100011011000010101011;
		correct = 32'b00110100100100001001000100111010;
		#400 //1.1956896e-26 * 4.4403608e-20 = 2.6927756e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011010110010010100000101111010;
		b = 32'b10010100011101110111101110010001;
		correct = 32'b11000101110100000010111010100001;
		#400 //8.3237435e-23 * -1.2494682e-26 = -6661.8286
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010110110010111101001011000001;
		b = 32'b10000101011000010011001001100110;
		correct = 32'b11010000111001111011001111101101;
		#400 //3.2929423e-25 * -1.0588706e-35 = -31098628000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010010011101010010110100110;
		b = 32'b00000110111001010111110010000101;
		correct = 32'b11110010111001101000010110011101;
		#400 //-0.000788296 * 8.632319e-35 = -9.1319143e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101010110111101111011011000111;
		b = 32'b11001011110100111000111011011011;
		correct = 32'b10011110100001101110011010101000;
		#400 //3.9606358e-13 * -27729334.0 = -1.4283199e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100101110010101001000001011111;
		b = 32'b01101001111111111110000000110010;
		correct = 32'b10111011010010101010100110001101;
		#400 //-1.1957265e+23 * 3.8666852e+25 = -0.0030923814
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101011100001110001110011000110;
		b = 32'b10101000110101111001001101101101;
		correct = 32'b01000010001000000111001011000001;
		#400 //-9.600313e-13 * -2.393373e-14 = 40.112064
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111111011011011000000110101101;
		b = 32'b10111010000000011110000101110101;
		correct = 32'b01000100111010100001000101000010;
		#400 //-0.92775995 * -0.0004954555 = 1872.5393
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010100000010011110110111100100;
		b = 32'b01101101010010001011101000111110;
		correct = 32'b10100110001011111110100011011010;
		#400 //-2369606600000.0 * 3.8826347e+27 = -6.1030894e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010100011100110110100000010111;
		b = 32'b11010000101111101110100011010100;
		correct = 32'b11000011001000110011001010110000;
		#400 //4181693600000.0 * -25623437000.0 = -163.198
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000011011001100110000111101110;
		b = 32'b00000111001110000000001100110011;
		correct = 32'b10111011101000000100000101010111;
		#400 //-6.7703343e-37 * 1.3843562e-34 = -0.0048906016
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000010011101001010101100111001;
		b = 32'b10011010101111111000111110100111;
		correct = 32'b10100111001000110111110001111010;
		#400 //1.7975427e-37 * -7.922783e-23 = -2.2688273e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101001011011011100000100001011;
		b = 32'b10101001000000011100010111011011;
		correct = 32'b10111111111010101000000110001011;
		#400 //5.279201e-14 * -2.8815366e-14 = -1.8320783
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000110000110001110011000101000;
		b = 32'b00101101011010100100101001100110;
		correct = 32'b01011000001001110001000100010010;
		#400 //9785.539 * 1.331788e-11 = 734767000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011100010101100101011100011101;
		b = 32'b11111001011111111000111000000000;
		correct = 32'b00100010010101101011011010111010;
		#400 //-2.413257e+17 * -8.293224e+34 = 2.9099143e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101110010011001100010111010110;
		b = 32'b01001111101011000010110000111001;
		correct = 32'b11011110000110000011110001110101;
		#400 //-1.5843528e+28 * 5777158700.0 = -2.7424429e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101101000000001100011000100011;
		b = 32'b10000111100110001100000011111000;
		correct = 32'b01100100110101111100111111101111;
		#400 //-7.319953e-12 * -2.2983835e-34 = 3.1848265e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111110001101011100100101110001;
		b = 32'b01101000101101111011001000100001;
		correct = 32'b11010100111111010101011011110110;
		#400 //-6.0409053e+37 * 6.939832e+24 = -8704685500000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101111011001011100111011110000;
		b = 32'b11011111010111010100110100010001;
		correct = 32'b00001111100001001110101110101101;
		#400 //-2.0900948e-10 * -1.594642e+19 = 1.3106984e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110101111100100100110100000101;
		b = 32'b01100011111000101000101001110001;
		correct = 32'b11010001100010001110011110011110;
		#400 //-6.1430566e+32 * 8.35788e+21 = -73500180000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111000001001010000000011011111;
		b = 32'b11111010001001000111110100101101;
		correct = 32'b10111101100000000110011001111011;
		#400 //1.3386666e+34 * -2.1351889e+35 = -0.062695466
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000011100111101001100111001;
		b = 32'b00110110010010101010101001001101;
		correct = 32'b10111001100110011111111011110010;
		#400 //-8.870305e-10 * 3.0199474e-06 = -0.00029372383
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000100001001010100111010001000;
		b = 32'b11010000011110111000011011101111;
		correct = 32'b00110011001010000011111100010101;
		#400 //-661.22705 * -16879697000.0 = 3.917292e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100111011011010110101010101010;
		b = 32'b00010011011000100000010110010111;
		correct = 32'b01010011100001100111001111111101;
		#400 //3.294818e-15 * 2.8527966e-27 = 1154943200000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111101001010000011111101100010;
		b = 32'b01010100111111111101110010010110;
		correct = 32'b00100111101010000101011010101100;
		#400 //0.04107607 * 8791340000000.0 = 4.6723337e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011010101001100101111110010100;
		b = 32'b10101000101001100000111101000011;
		correct = 32'b11110001100000000011110111101001;
		#400 //2.3414968e+16 * -1.8436321e-14 = -1.2700456e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100110011101001101110111000111;
		b = 32'b00000100110010010110010111010111;
		correct = 32'b11100001000110111010000001110011;
		#400 //-8.495507e-16 * 4.7348398e-36 = -1.7942543e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001100110100000100101110100011;
		b = 32'b01101100010110101110101011011001;
		correct = 32'b00011111111100111001010000101110;
		#400 //109206810.0 * 1.05861946e+27 = 1.03159646e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011100011110000111000100100101;
		b = 32'b01000110110111110111101001001010;
		correct = 32'b01010101000011100100110001110100;
		#400 //2.797208e+17 * 28605.145 = 9778688000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011001000010001011110101101010;
		b = 32'b10010001000010101000111110001010;
		correct = 32'b01000111011111001010001011001110;
		#400 //-7.069287e-24 * -1.0930512e-28 = 64674.805
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100111011111000100101011100;
		b = 32'b11101011011010010100101010100001;
		correct = 32'b10011001000000110110110100101101;
		#400 //1916.2925 * -2.8203214e+26 = -6.794589e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000101101001011010101111001100;
		b = 32'b00001001110110011011110010000011;
		correct = 32'b10111011010000101100100011111011;
		#400 //-1.5579634e-35 * 5.2418125e-33 = -0.0029721844
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101110011111000111011000010010;
		b = 32'b11010011100101101111111000111001;
		correct = 32'b01011010010101100000010001000110;
		#400 //-1.953324e+28 * -1297020500000.0 = 1.5060086e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111101111111000001001000001000;
		b = 32'b01001111010111010001001011000001;
		correct = 32'b11101110000100011111001001111010;
		#400 //-4.1882385e+37 * 3708993800.0 = -1.1292116e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011010110011100100001101101110;
		b = 32'b11101101010101100100101110001111;
		correct = 32'b10101100111101100110011110111000;
		#400 //2.9028992e+16 * -4.145071e+27 = -7.0032556e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011011010010100111010010101111;
		b = 32'b00001010100100100000010010001000;
		correct = 32'b01010000001100010111100101010110;
		#400 //1.6746751e-22 * 1.4060993e-32 = 11910076000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001111101111100101000000101000;
		b = 32'b00100001101010010101110101011011;
		correct = 32'b01101101100011111101010100000101;
		#400 //6385848300.0 * 1.1476596e-18 = 5.564235e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100100000011000100000100111111;
		b = 32'b11010110010000111000110000100110;
		correct = 32'b00001101001101111001110100101110;
		#400 //-3.0412926e-17 * -53751675000000.0 = 5.6580427e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000000010001011101010101000111;
		b = 32'b01011010001011010000011110111000;
		correct = 32'b00100101100100100101100100011111;
		#400 //3.0911424 * 1.2175914e+16 = 2.5387354e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011011000000111111111111110001;
		b = 32'b01001001111101111100110010100001;
		correct = 32'b10010000100010000101111001000000;
		#400 //-1.0918765e-22 * 2029972.1 = -5.3787757e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110011100001101000101100110100;
		b = 32'b11011101010100110000000010001011;
		correct = 32'b01010101101000110011110001111101;
		#400 //-2.131931e+31 * -9.502691e+17 = 22435024000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010010000100011101100000011010;
		b = 32'b00101010111000111010011110011000;
		correct = 32'b10100110101001000000000011010100;
		#400 //-4.60203e-28 * 4.0439592e-13 = -1.138001e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111110111110011111001010010101;
		b = 32'b11011000100000100001000111000101;
		correct = 32'b01100101111101011111100010001101;
		#400 //-1.6611866e+38 * -1144102600000000.0 = 1.4519559e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000111000101110011100101111101;
		b = 32'b10111001100111110011110111001101;
		correct = 32'b00001100111100110001110010101000;
		#400 //-1.1376872e-34 * -0.00030372888 = 3.7457325e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000110111000011101111110010111;
		b = 32'b10000001010111101111001101000100;
		correct = 32'b11000101000000011010110110100001;
		#400 //8.496413e-35 * -4.0949495e-38 = -2074.8518
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101001011011101001001001110101;
		b = 32'b10101110001010001100111101111111;
		correct = 32'b10111010101101001110010101111111;
		#400 //5.2973647e-14 * -3.838307e-11 = -0.0013801305
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100101101001101010111100100;
		b = 32'b10001010000001000100011001011100;
		correct = 32'b11111010001011101111110111000101;
		#400 //1446.6841 * -6.368802e-33 = -2.2715168e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011000010100010101011000110011;
		b = 32'b10110010010000110001000011110011;
		correct = 32'b10100101100010010101110100111000;
		#400 //2.7056136e-24 * -1.1354348e-08 = -2.382888e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101000110011010100100000110111;
		b = 32'b10010001100110100110001100100000;
		correct = 32'b01010110101010100011001000110111;
		#400 //-2.279089e-14 * -2.4358006e-28 = 93566320000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011101111010100000001101010010;
		b = 32'b01001000000100100000001000001111;
		correct = 32'b01010101010011010010011010011000;
		#400 //2.1078014e+18 * 149512.23 = 14097853000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001101001101010101100001110111;
		b = 32'b11001000100001101111100010100000;
		correct = 32'b11000100001010111111101010101010;
		#400 //190154610.0 * -276421.0 = -687.9166
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000110001011011111011101001001;
		b = 32'b00001101111100110101101111101010;
		correct = 32'b10110111101101110000000010011100;
		#400 //-3.271936e-35 * 1.4998159e-30 = -2.1815584e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111001100100001111101010010010;
		b = 32'b00100011001100001001111001000111;
		correct = 32'b11010101110100100010001111011010;
		#400 //-0.0002765251 * 9.574496e-18 = -28881428000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010011101101100011101010111101;
		b = 32'b10011001011010000000100001010100;
		correct = 32'b01111001110010010000110101110110;
		#400 //-1565339000000.0 * -1.1995801e-23 = 1.3049059e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010110111100110100011001100111;
		b = 32'b01011110011010100110111010111001;
		correct = 32'b00111000000001001101001111111000;
		#400 //133741850000000.0 * 4.2231607e+18 = 3.1668664e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001110001000010001010101100011;
		b = 32'b01001001110000111000100101011110;
		correct = 32'b10000011110100101110010010111001;
		#400 //-1.985508e-30 * 1601835.8 = -1.2395203e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010101101110101011010000111000;
		b = 32'b10100100100011100010011001010001;
		correct = 32'b11110000101010000001111010001101;
		#400 //25660400000000.0 * -6.1647594e-17 = -4.1624332e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111111100010010111110001010101;
		b = 32'b11011001001100111000001110010101;
		correct = 32'b00100101110001000001000010000111;
		#400 //-1.0741068 * -3158043600000000.0 = 3.401178e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101101101110111000010010001011;
		b = 32'b10110001100001001111111110110000;
		correct = 32'b01111011101101000111100001001001;
		#400 //-7.2542414e+27 * -3.870774e-09 = 1.8741062e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111111010001001011011010110000;
		b = 32'b00001111000001010001101100011001;
		correct = 32'b11101111101111010010101011110110;
		#400 //-0.7684126 * 6.562625e-30 = -1.1708921e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100110101111100111011000110010;
		b = 32'b01111111110110100011001000010101;
		correct = 32'b01111111110110100011001000010101;
		#400 //-1.3215935e-15 * nan = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011101001001111011100100000100;
		b = 32'b10001001010001100000111111011111;
		correct = 32'b11010011010110001100100100100110;
		#400 //2.2197917e-21 * -2.3840846e-33 = -931087650000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100100100010010111010111111001;
		b = 32'b11001011011010111101110111111101;
		correct = 32'b11011000100101010011000110101101;
		#400 //2.0285638e+22 * -15457789.0 = -1312324700000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111001000101101000010101010001;
		b = 32'b11011101101011000101001001100111;
		correct = 32'b00011010110111111001110011001001;
		#400 //-0.00014354779 * -1.5521375e+18 = 9.248394e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111101101001101011011111010010;
		b = 32'b11111010100110011001010100101111;
		correct = 32'b11000010100010101111001010000011;
		#400 //2.7700787e+37 * -3.987236e+35 = -69.473656
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111100110110111111101100110111;
		b = 32'b11111011000010111101011010011101;
		correct = 32'b10000001010010010101101110111001;
		#400 //0.026853187 * -7.260821e+35 = -3.6983677e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101010001001110010101000011111;
		b = 32'b10001101000011001011110101111011;
		correct = 32'b01011100100110000000100001001010;
		#400 //-1.4847193e-13 * -4.336891e-31 = 3.423465e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010011101011101001011001000101;
		b = 32'b01011001101101011001010000111110;
		correct = 32'b10111001011101100010010001100110;
		#400 //-1499690800000.0 * 6388745600000000.0 = -0.00023473948
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000010011011001100010110000011;
		b = 32'b00011001100000000111111010001100;
		correct = 32'b11101000011010111101110001010100;
		#400 //-59.192883 * 1.3286002e-23 = -4.4552818e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110001111101001110111000111000;
		b = 32'b11001110011001001111011101111001;
		correct = 32'b11100011000010001110110010100001;
		#400 //2.4256746e+30 * -960355900.0 = -2.525808e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111110000101001101111011111;
		b = 32'b10001100111011001101000100100011;
		correct = 32'b01101010010100100101111101111000;
		#400 //-2.3199185e-05 * -3.6487427e-31 = 6.3581315e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001101010011011110111010101000;
		b = 32'b00010110111010000011001111110000;
		correct = 32'b00110101111000110000100101111100;
		#400 //6.3457774e-31 * 3.7514399e-25 = 1.6915578e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101101110111100011110001110010;
		b = 32'b11101000001010110001100010010000;
		correct = 32'b01000101001001100100001001000111;
		#400 //-8.597343e+27 * -3.231911e+24 = 2660.1423
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001011101000101100011011101101;
		b = 32'b10100010101101011001100101110110;
		correct = 32'b10101000011001010111011101010101;
		#400 //6.269944e-32 * -4.922263e-18 = -1.273793e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010010001100010100110101001100;
		b = 32'b10000101111010110111101010001001;
		correct = 32'b01001011110000001100000011011011;
		#400 //-5.594663e-28 * -2.2144306e-35 = 25264566.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010011011101000111101001110011;
		b = 32'b01000101011001010100010110100111;
		correct = 32'b11001101100010000111110101001110;
		#400 //-1050026400000.0 * 3668.3533 = -286239170.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110110011101010010000101000110;
		b = 32'b00100111011000100001111010000101;
		correct = 32'b01001110100010101100001011110000;
		#400 //3.6527213e-06 * 3.1380345e-15 = 1164015600.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110111001110000111101101110110;
		b = 32'b11000110010010000000110000011011;
		correct = 32'b01110000011011000001010011011100;
		#400 //-3.741745e+33 * -12803.026 = 2.9225472e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101111100101111000100100111011;
		b = 32'b11011001101001010000011011110110;
		correct = 32'b11010101011010110001001001011110;
		#400 //9.379628e+28 * -5806378000000000.0 = -16154007000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011111011010100100000110110110;
		b = 32'b01001000011001101101100100101010;
		correct = 32'b10010110100000011110001111001111;
		#400 //-4.9605782e-20 * 236388.66 = -2.0984841e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100001100010101000111100110111;
		b = 32'b01000111111100100100001010001001;
		correct = 32'b10011001000100100110101100000011;
		#400 //-9.389152e-19 * 124037.07 = -7.569634e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101100001000001101000001101001;
		b = 32'b00111111001101001110101100000111;
		correct = 32'b01101100011000111000110110000011;
		#400 //7.776493e+26 * 0.70671123 = 1.1003777e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110110110001110111010100010010;
		b = 32'b11001001100000000010100100101111;
		correct = 32'b11101100110001110011010011111010;
		#400 //2.0227374e+33 * -1049893.9 = -1.9266113e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001101011110001000001110011000;
		b = 32'b11000101000111101011111010001001;
		correct = 32'b11000111110010000110001001000111;
		#400 //260585860.0 * -2539.9084 = -102596.555
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001100011001101000001010101001;
		b = 32'b10100100111011111000000000101001;
		correct = 32'b11100110111101100110001111110011;
		#400 //60426916.0 * -1.0386684e-16 = -5.8177295e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111100110000110011001101001010;
		b = 32'b11100001111101100101010000111100;
		correct = 32'b01011010010010101101110100101110;
		#400 //-8.108305e+36 * -5.679961e+20 = 1.4275284e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001011001001101001001110110110;
		b = 32'b00110001100011011111100010001010;
		correct = 32'b10011001000101100010111101001011;
		#400 //-3.2081562e-32 * 4.1318957e-09 = -7.764369e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111011111011001100001101001111;
		b = 32'b01101111110110001100011001111000;
		correct = 32'b10001011100010111100110101011011;
		#400 //-0.007225431 * 1.3417739e+29 = -5.3849837e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111110011001111010111100011;
		b = 32'b11001011011000111100010111010010;
		correct = 32'b10111011111001100101110001010111;
		#400 //104939.77 * -14927314.0 = -0.0070300507
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001111100010100101100011001011;
		b = 32'b00100000110010010110010100100000;
		correct = 32'b00101110001011111101101101111011;
		#400 //1.3642052e-29 * 3.4117643e-19 = 3.998533e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001111001000110111110100001101;
		b = 32'b11111010010100011010101010010110;
		correct = 32'b00010100010001111001111000001110;
		#400 //-2742881500.0 * -2.7216248e+35 = 1.0078103e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111101100010100101110011100000;
		b = 32'b00010011010001001010111000111011;
		correct = 32'b11101001101101000001011111101001;
		#400 //-0.06755996 * 2.482458e-27 = -2.7214945e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000111111000010100000011100000;
		b = 32'b00001110001101100101100010111111;
		correct = 32'b10111001000111100001111001101010;
		#400 //-3.3892367e-34 * 2.2475962e-30 = -0.00015079384
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011001011101010100011110110100;
		b = 32'b10110111100111100000100001010001;
		correct = 32'b01100001010001101010101011000101;
		#400 //-4315013000000000.0 * -1.883894e-05 = 2.2904754e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101111001110111111001101110001;
		b = 32'b11000001000101001000101100100011;
		correct = 32'b01101101101000011111010100011001;
		#400 //-5.8168e+28 * -9.283969 = 6.265424e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010100110010111000101011011001;
		b = 32'b10000000111011111111110111100101;
		correct = 32'b11010011010110010001111010001011;
		#400 //2.0552528e-26 * -2.2039764e-38 = -932520300000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100001100010000110000100110101;
		b = 32'b11100001111101100000100001100110;
		correct = 32'b00111111000011011110011110011001;
		#400 //-3.144702e+20 * -5.6731303e+20 = 0.55431515
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101010111101100001100011100101;
		b = 32'b11000100101110100010010100101110;
		correct = 32'b00100101101010010011100110100001;
		#400 //-4.3715652e-13 * -1489.1619 = 2.9355878e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001000101001101110000100001011;
		b = 32'b01000111111000100101000000110111;
		correct = 32'b11000000001111001100010011111010;
		#400 //-341768.34 * 115872.43 = -2.9495225
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101011001010110100001100111011;
		b = 32'b10110001100100111001100010001001;
		correct = 32'b11111001000101001000011001001101;
		#400 //2.070438e+26 * -4.2956043e-09 = -4.819899e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110100101100000010010010011001;
		b = 32'b01110011101010101100011010000001;
		correct = 32'b11000000100001000000010111101010;
		#400 //-1.1164386e+32 * 2.7060443e+31 = -4.125722
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000011000011100010000010100101;
		b = 32'b00111100010010111101010011100011;
		correct = 32'b11000110001100101000000011100011;
		#400 //-142.12752 * 0.012440893 = -11424.222
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101001110111110011000011000111;
		b = 32'b11000011001010111011011000111110;
		correct = 32'b10100110001001100101111110111101;
		#400 //9.911651e-14 * -171.71188 = -5.772257e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111101011111011101001001011010;
		b = 32'b01001001100111101011000001110000;
		correct = 32'b10110011010011001011110000010000;
		#400 //-0.061968185 * 1299982.0 = -4.7668493e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111101100011110001100101101011;
		b = 32'b11011000011000000101011000001101;
		correct = 32'b01100100101000110100110000001000;
		#400 //-2.3776448e+37 * -986640760000000.0 = 2.4098383e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101001000001010110101011001101;
		b = 32'b01000011101100101100110001000110;
		correct = 32'b01100100101111110000011001001010;
		#400 //1.0080718e+25 * 357.5959 = 2.819025e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000001100001110001100100010111;
		b = 32'b00001011010100100000001110010100;
		correct = 32'b10110101101001001010111000010001;
		#400 //-4.962717e-38 * 4.044722e-32 = -1.2269612e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101011111000010101010000110011;
		b = 32'b11000001110100100001101101011110;
		correct = 32'b10101001100010010100011000000001;
		#400 //1.6010582e-12 * -26.263363 = -6.096166e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010000001110001111000010110010;
		b = 32'b01100101110000100001010000011000;
		correct = 32'b10101001111100111111001000110101;
		#400 //-12411128000.0 * 1.1456372e+23 = -1.0833384e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101100001001000110100111110100;
		b = 32'b00001110111100000111100110100110;
		correct = 32'b01011100101011110000011100111100;
		#400 //2.3364618e-12 * 5.928171e-30 = 3.941286e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100010000011000101100011101011;
		b = 32'b11000100110101000111001001110010;
		correct = 32'b00011100101010010001111010010001;
		#400 //-1.902061e-18 * -1699.5764 = 1.1191383e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100001011100011001111010100011;
		b = 32'b00100100111011010001000100101011;
		correct = 32'b11111100000000100111010101000110;
		#400 //-2.7856852e+20 * 1.0281145e-16 = -2.7095087e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101110110011010101000100101010;
		b = 32'b01010101010100100001111111010101;
		correct = 32'b11011000111110100010010010100101;
		#400 //-3.1771274e+28 * 14439635000000.0 = -2200282400000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000011110100111011010001010100;
		b = 32'b00000100111101011010100110110101;
		correct = 32'b11111110010111001001110011010001;
		#400 //-423.4088 * 5.7755074e-36 = -7.33111e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111100000111000110010111111111;
		b = 32'b01111000111000001100010100011100;
		correct = 32'b11000010101100100010000011110111;
		#400 //-3.248268e+36 * 3.647101e+34 = -89.064384
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000111010000001100001100011000;
		b = 32'b01101111100111010111101101101001;
		correct = 32'b10010111000111001010110011011111;
		#400 //-49347.094 * 9.747668e+28 = -5.0624513e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111100110010111001011110111;
		b = 32'b10111111100111011100100001000001;
		correct = 32'b00110111011110001111100000110001;
		#400 //-1.8292556e-05 * -1.2326738 = 1.48397385e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000110010010100001000110100010;
		b = 32'b10100100111011010100100111011101;
		correct = 32'b01100000110110100000000011001011;
		#400 //-12932.408 * -1.02907495e-16 = 1.2567023e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111011010101110001100010111;
		b = 32'b00111011010101100011001001000111;
		correct = 32'b01001011100011000101110101001000;
		#400 //60131.09 * 0.0032683776 = 18397840.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110110111010100101010000010001;
		b = 32'b11001100000011110000011110111110;
		correct = 32'b11101010010100011011010001000010;
		#400 //2.3763721e+33 * -37494520.0 = -6.3379185e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001000100111110101000011101111;
		b = 32'b10010100001111110110010011100110;
		correct = 32'b00110011110101010001100000001110;
		#400 //-9.588492e-34 * -9.6629344e-27 = 9.922961e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100001000001101100100001110010;
		b = 32'b11010111100011111011101110000000;
		correct = 32'b01001000111100000000111101101110;
		#400 //-1.553942e+20 * -316070940000000.0 = 491643.44
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110010101000001101101110110000;
		b = 32'b11100100001000001110010000100011;
		correct = 32'b01001101111111111111001010001110;
		#400 //-6.372248e+30 * -1.1871672e+22 = 536760770.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101001110001100010011111001000;
		b = 32'b01010101001101110010111010011000;
		correct = 32'b00010100000010100111011001111001;
		#400 //8.799867e-14 * 12588172000000.0 = 6.990584e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101001110101000001010001101111;
		b = 32'b11100001110110010000000110011010;
		correct = 32'b00000111011110100011000000110111;
		#400 //-9.418236e-14 * -5.0038236e+20 = 1.8822079e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000001110011101111001001001001;
		b = 32'b00011100110000001111001111111011;
		correct = 32'b01100100100010010100100001101000;
		#400 //25.868303 * 1.2768562e-21 = 2.025937e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000001100101100001111111111010;
		b = 32'b11011000010111010100111000101111;
		correct = 32'b10101000101011011010100100001101;
		#400 //18.765614 * -973311460000000.0 = -1.9280172e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110011000101101111000010011100;
		b = 32'b01000111111010110101001011011101;
		correct = 32'b11101010101001000011001110110011;
		#400 //-1.1958689e+31 * 120485.73 = -9.925399e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101001101111100010111110001010;
		b = 32'b00100011100101110011110011010111;
		correct = 32'b01000101101000001111011010110100;
		#400 //8.445942e-14 * 1.639722e-17 = 5150.838
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011001110011000101010100000000;
		b = 32'b10101000110000101110101000110100;
		correct = 32'b11110000100001100010111100101010;
		#400 //7189294000000000.0 * -2.1639896e-14 = -3.3222407e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010110011101100001100100010101;
		b = 32'b00101100110000111101110110011011;
		correct = 32'b01101001001000001101001111001001;
		#400 //67646897000000.0 * 5.5668365e-12 = 1.2151766e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101000011101111010001010010101;
		b = 32'b01011101110100011000000000101111;
		correct = 32'b01001010000101110100110010011000;
		#400 //4.6776945e+24 * 1.8870147e+18 = 2478886.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100010110111111100111000010000;
		b = 32'b10110000010011110011111101011011;
		correct = 32'b00110010000010100011100111101000;
		#400 //-6.066245e-18 * -7.5396195e-10 = 8.045824e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010000100001101110101010001011;
		b = 32'b10010000001101001101001101001010;
		correct = 32'b10111111101111110000000101000111;
		#400 //5.321505e-29 * -3.5661512e-29 = -1.4922265
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111000111011110011001011100001;
		b = 32'b11010111010100010000110111000101;
		correct = 32'b11100001000100100111010100001101;
		#400 //3.8812216e+34 * -229857070000000.0 = -1.6885369e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101001001101000110111110001011;
		b = 32'b10100111110101011011010111111000;
		correct = 32'b11000000110110000010001111110010;
		#400 //4.0064777e-14 * -5.9316667e-15 = -6.754388
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100001101100110010010101010000;
		b = 32'b10100100000100000001010110001101;
		correct = 32'b10111101000111110010010111001011;
		#400 //1.2139388e-18 * -3.1243277e-17 = -0.0388544
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011000100011011101101001010000;
		b = 32'b00101100010001000000001010101111;
		correct = 32'b01101011101110010100010001100111;
		#400 //1247750300000000.0 * 2.7854765e-12 = 4.479486e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111011110000100001011111110011;
		b = 32'b00111101001010100101000110011000;
		correct = 32'b11111110000100011101111000011000;
		#400 //-2.0155827e+36 * 0.04158172 = -4.847281e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011101100010010000000010000110;
		b = 32'b10010000110100000110100001100001;
		correct = 32'b01001100001010000100100110111011;
		#400 //-3.626414e-21 * -8.2202355e-29 = 44115692.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010111011100101111110101001111;
		b = 32'b11001011001101000011000001111100;
		correct = 32'b00001011101011001001110001100100;
		#400 //-7.851414e-25 * -11808892.0 = 6.64873e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111101011011011111100000000110;
		b = 32'b01011111001010111000101111000000;
		correct = 32'b01011101101100011000111111010111;
		#400 //1.9769678e+37 * 1.2361185e+19 = 1.5993352e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001000110110101111111010111100;
		b = 32'b11000001111111010101011101101001;
		correct = 32'b00000110010111010100101100001110;
		#400 //-1.31802855e-33 * -31.66768 = 4.1620622e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110000110111011010100111011;
		b = 32'b00110000110001000101011001101100;
		correct = 32'b01001100110010110000011000100001;
		#400 //0.15205853 * 1.428544e-09 = 106443016.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100111011100011011001111100101;
		b = 32'b00011101000011000110111010000000;
		correct = 32'b01001001110111000100111001011101;
		#400 //3.354299e-15 * 1.8585973e-21 = 1804747.6
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000011110111100011101010010110;
		b = 32'b11100011101101000101011110110000;
		correct = 32'b00011111100111011011101010110001;
		#400 //-444.4577 * -6.653465e+21 = 6.680094e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000010100101011100011110011000;
		b = 32'b11111001110101100100011000000010;
		correct = 32'b10001000001100101111001001101110;
		#400 //74.88983 * -1.3907143e+35 = -5.38499e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111101010110100110111111111011;
		b = 32'b01000100010111010111110011010110;
		correct = 32'b01111000011111000111100101111001;
		#400 //1.8147071e+37 * 885.95056 = 2.0483165e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010010111111101110010110011;
		b = 32'b01100110010010001000000110100010;
		correct = 32'b10010011100011101110100011110000;
		#400 //-0.00085396616 * 2.3671615e+23 = -3.6075534e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101100110000111111101111101010;
		b = 32'b10000011000000101001011110101100;
		correct = 32'b01101001010000000001011111101100;
		#400 //-5.5702014e-12 * -3.8377677e-37 = 1.451417e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010101101010100110011111111010;
		b = 32'b10101110101111011001111001010011;
		correct = 32'b10100110011001100000111111010111;
		#400 //6.88265e-26 * -8.622849e-11 = -7.9818747e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000101011001100000101001100100;
		b = 32'b01110111010001101000101011100001;
		correct = 32'b10001101100101000100111010001000;
		#400 //-3680.6494 * 4.0269202e+33 = -9.14011e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101111111110010011011100100101;
		b = 32'b11110100000100100101011001010101;
		correct = 32'b00111011010110011111110010011001;
		#400 //-1.5425687e+29 * -4.637612e+31 = 0.0033262132
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011010010010010010000000001101;
		b = 32'b11010110110001011100100110101101;
		correct = 32'b01000011000000100010100011101010;
		#400 //-1.4152928e+16 * -108734990000000.0 = 130.15982
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110011111100000101111100011110;
		b = 32'b10111101101111100001011100111101;
		correct = 32'b10110101101000011101101101110001;
		#400 //1.11931726e-07 * -0.09281776 = -1.2059301e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101001000110001100110101001101;
		b = 32'b00001111101101011110110101010001;
		correct = 32'b01011000110101110000010000110110;
		#400 //3.392885e-14 * 1.7939389e-29 = 1891304700000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100010011000101100100101100111;
		b = 32'b11000100000000000110011000110001;
		correct = 32'b01011101111000100001010011101000;
		#400 //-1.0458692e+21 * -513.59674 = 2.0363626e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010000010010010011110110001111;
		b = 32'b00111101111010100001001001101110;
		correct = 32'b01010001110111000001011111000001;
		#400 //13505019000.0 * 0.114292964 = 118161420000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000110110001100011101000010010;
		b = 32'b10001001110001000111100101101000;
		correct = 32'b00111100100000010010010001001100;
		#400 //-7.456465e-35 * -4.7299454e-33 = 0.015764378
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111001111010100010000010110001;
		b = 32'b00010101001111100100001101100011;
		correct = 32'b01100100000111011000001010001010;
		#400 //0.00044656315 * 3.8423353e-26 = 1.1622181e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000100011110001111000100011100;
		b = 32'b00100001010101011001101010110110;
		correct = 32'b00100010100101010010110011110100;
		#400 //2.9262972e-36 * 7.2371965e-19 = 4.0434127e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110101011110001001100110110000;
		b = 32'b10000010000001111001111111001010;
		correct = 32'b01110010111010101010000000001010;
		#400 //-9.2610844e-07 * -9.964091e-38 = 9.29446e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110111111001001110011010001110;
		b = 32'b00101100110101011111111101110111;
		correct = 32'b01001010100010001110100111110010;
		#400 //2.7287078e-05 * 6.0821864e-12 = 4486393.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101000111110001101100011101000;
		b = 32'b01001010010110111101100111001110;
		correct = 32'b01011110000100001110000111010100;
		#400 //9.401185e+24 * 3602035.5 = 2.6099646e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011010001110100101101000110000;
		b = 32'b11110100000001111100101110000100;
		correct = 32'b10100101101011111010011110111011;
		#400 //1.3113377e+16 * -4.303515e+31 = -3.047132e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000001010100000111101110101010;
		b = 32'b00001100011101100011100001000011;
		correct = 32'b10110100010110001100001110101011;
		#400 //-3.829229e-38 * 1.8968081e-31 = -2.0187751e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011101010010011110000001010101;
		b = 32'b10000011000110111011111001101010;
		correct = 32'b01011001101001011110101000100001;
		#400 //-2.6718105e-21 * -4.576899e-37 = 5837600000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000001010001000101110010010111;
		b = 32'b11110000101001111010010111110111;
		correct = 32'b00010000000101011110110000111010;
		#400 //-12.272605 * -4.150771e+29 = 2.956705e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010100011110011000010100100100;
		b = 32'b00100110101010001111110101001001;
		correct = 32'b00101101001111001111111101011011;
		#400 //1.2597545e-26 * 1.1725995e-15 = 1.0743263e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010010110011011100110101110011;
		b = 32'b11110000100001010110011111101001;
		correct = 32'b10100001110001010111011010000101;
		#400 //441957580000.0 * -3.30297e+29 = -1.3380611e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100001011000001111111101111001;
		b = 32'b10100001101001110011101000000111;
		correct = 32'b01111111001011000011100001000010;
		#400 //-2.5940496e+20 * -1.133172e-18 = 2.2891932e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011100010100100001101110010110;
		b = 32'b11011000010000111010001111100001;
		correct = 32'b01000011100010010111011100110010;
		#400 //-2.365603e+17 * -860434500000000.0 = 274.9312
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010011010100001010110111101010;
		b = 32'b00011011001100011001111100010010;
		correct = 32'b11110111100101100110000110100110;
		#400 //-896271000000.0 * 1.4692495e-22 = -6.100196e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100000001111101000011001100000;
		b = 32'b10000000010011001110000001010000;
		correct = 32'b01011111100111101001110100000100;
		#400 //-1.6138087e-19 * -7.059966e-39 = 2.2858592e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000100010110011111100101011011;
		b = 32'b10100000101101000100011000111000;
		correct = 32'b10100011000110101100010010010111;
		#400 //2.5622726e-36 * -3.0539653e-19 = -8.389986e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110100111011000101100100101101;
		b = 32'b00010111100010011011100110011000;
		correct = 32'b01011100110110111010100011010000;
		#400 //4.402331e-07 * 8.900268e-25 = 4.9462905e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001010100101001101001100101001;
		b = 32'b00010011111100011100011010001011;
		correct = 32'b01110110000111011001010010101000;
		#400 //4876692.5 * 6.103273e-27 = 7.99029e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100010110101011111000001111111;
		b = 32'b01111101011000000100010001100001;
		correct = 32'b00100100111101000011011000000101;
		#400 //1.973243e+21 * 1.8631382e+37 = 1.05909645e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111100000101011110001100001001;
		b = 32'b10111111011001110111010000010010;
		correct = 32'b10111100001001011100100001110010;
		#400 //0.009148368 * -0.90411484 = -0.010118591
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000101011000010011100101010;
		b = 32'b01000111011000111011011111101110;
		correct = 32'b10101000110000011000100010010110;
		#400 //-1.2525778e-09 * 58295.93 = -2.1486539e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000100011010001010000111101110;
		b = 32'b00010100110000110100011110111100;
		correct = 32'b11101111000110000111101110110111;
		#400 //-930.53015 * 1.9718262e-26 = -4.7191284e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000111111011110000101011011010;
		b = 32'b10101100001100000001111101011100;
		correct = 32'b10011011001011011011101001100100;
		#400 //3.5967101e-34 * -2.5028512e-12 = -1.4370451e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100000011011011101011101010001;
		b = 32'b01010101001001010000010100010100;
		correct = 32'b10001010101110000111110000011111;
		#400 //-2.0145923e-19 * 11340077000000.0 = -1.7765245e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010101100110111011010100101001;
		b = 32'b10110000000110011101100010100100;
		correct = 32'b10100101000000011000110001110111;
		#400 //6.288982e-26 * -5.596894e-10 = -1.1236558e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110010010100000100010000110000;
		b = 32'b01010101110110011111011001111111;
		correct = 32'b10011011111101001001110010000000;
		#400 //-1.21226975e-08 * 29956590000000.0 = -4.046755e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100010000001010111101010000011;
		b = 32'b01011000100100110010010001110000;
		correct = 32'b11001000111010000011101001000100;
		#400 //-6.155612e+20 * 1294277700000000.0 = -475602.12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110111101101001001111001001111;
		b = 32'b11100000101000100010011010111011;
		correct = 32'b10010110100011101001001111100011;
		#400 //2.153139e-05 * -9.3473855e+19 = -2.3034667e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100100001101111111011000010011;
		b = 32'b11011110111110100101100111110000;
		correct = 32'b00000100101111000001110010101001;
		#400 //-3.9890232e-17 * -9.019857e+18 = 4.4224908e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101101001100000100000111110000;
		b = 32'b10100111011110100100111111100010;
		correct = 32'b11000101001101000100001101000100;
		#400 //1.0019083e-11 * -3.4737774e-15 = -2884.204
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000100011111100011001111101110;
		b = 32'b00100011100010000101001010010110;
		correct = 32'b00100000011011101010111011111110;
		#400 //2.9881401e-36 * 1.4780126e-17 = 2.0217284e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100011001110110001011110100111;
		b = 32'b00110011010010000100010001110100;
		correct = 32'b11101111011011110010100010010100;
		#400 //-3.4512455e+21 * 4.6628386e-08 = -7.4015973e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110011010110101011101101110011;
		b = 32'b11010000011101100000111100111001;
		correct = 32'b10100010011000111001000110011011;
		#400 //5.0927564e-08 * -16512771000.0 = -3.084132e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110100101010001000010011001111;
		b = 32'b11100101110111011110101101000101;
		correct = 32'b01001110010000100110011000011101;
		#400 //-1.0681147e+32 * -1.3099787e+23 = 815368000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010001001110101010100000100110;
		b = 32'b10000010011011101101110000001000;
		correct = 32'b01001110010010000000110100100001;
		#400 //-1.4724628e-28 * -1.7548624e-37 = 839075900.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011000111100001001001000000100;
		b = 32'b00101000010100101010111011000000;
		correct = 32'b11110000000100100010100010000101;
		#400 //-2116079400000000.0 * 1.1695235e-14 = -1.8093519e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011000110011010001100010001101;
		b = 32'b11001110000101101111100011111000;
		correct = 32'b01001010001011011110001101000100;
		#400 //-1804042600000000.0 * -633224700.0 = 2848977.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110001001100001100111100000011;
		b = 32'b00100011000101111011001001000111;
		correct = 32'b11001101100101010011000010000010;
		#400 //-2.5729043e-09 * 8.223478e-18 = -312873020.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101111100011111000010101100100;
		b = 32'b10010001011111110110110011011110;
		correct = 32'b11011101100011111101100000010000;
		#400 //2.6106328e-10 * -2.01495e-28 = -1.2956315e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010000110100111011011111001101;
		b = 32'b00010110110100001101111111110011;
		correct = 32'b00111001100000011011111000001000;
		#400 //8.3508015e-29 * 3.3745544e-25 = 0.00024746382
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010011101110010110001111001110;
		b = 32'b00110110110000111010100101111001;
		correct = 32'b10011100011100101000111101100110;
		#400 //-4.679898e-27 * 5.831182e-06 = -8.025642e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010110010010111110111100000111;
		b = 32'b11100011110011100101000100011001;
		correct = 32'b10110001111111010000101100000101;
		#400 //56056870000000.0 * -7.611746e+21 = -7.364522e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101111001100011011010001001100;
		b = 32'b10111000000000111011111110000111;
		correct = 32'b10110110101011001010011000010010;
		#400 //1.616211e-10 * -3.1411208e-05 = -5.1453326e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010001000100011011101000111000;
		b = 32'b00000011010100111000010110000101;
		correct = 32'b11001101001100000101111011101010;
		#400 //-1.1495866e-28 * 6.21606e-37 = -184938140.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011100001111100111000101110010;
		b = 32'b10111001001111100010001111100011;
		correct = 32'b01100010100000000011010000110110;
		#400 //-2.1441992e+17 * -0.00018133181 = 1.1824727e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100011101000100011100110000010;
		b = 32'b00011101110110111011010010001101;
		correct = 32'b01000101001111010000011000010010;
		#400 //1.758843e-17 * 5.8155502e-21 = 3024.3794
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100110110100100001011011111100;
		b = 32'b00001000101100000011011100110101;
		correct = 32'b11011101100110001001101100000111;
		#400 //-1.4577907e-15 * 1.0605594e-33 = -1.3745488e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001110011110101101001101111001;
		b = 32'b01101101001101100111100101110100;
		correct = 32'b10100000101011111111001001001110;
		#400 //-1052040770.0 * 3.5295687e+27 = -2.9806497e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011101100111101101010110000111;
		b = 32'b00110011111011111111111101111111;
		correct = 32'b11101001001010010110110010100111;
		#400 //-1.4306503e+18 * 1.1175779e-07 = -1.2801347e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010010011001001101111111110000;
		b = 32'b01110111111010110101010011110001;
		correct = 32'b00011001111110001111100111010010;
		#400 //245752400000.0 * 9.546192e+33 = 2.57435e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110011001111110100000000111111;
		b = 32'b00101001101000111101000111100100;
		correct = 32'b01001001000101010110111011100100;
		#400 //4.4529084e-08 * 7.2750643e-14 = 612078.25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001100001111010011110010111011;
		b = 32'b10110100011000100011011011001110;
		correct = 32'b01010111010101100010011110000100;
		#400 //-49607404.0 * -2.1067828e-07 = 235465200000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111001100011011100000011100000;
		b = 32'b00110101011111011101001001100011;
		correct = 32'b01000011100011101111100001001010;
		#400 //0.0002703732 * 9.4556e-07 = 285.93976
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011000100010100001010001001000;
		b = 32'b11001100101100100110100001111001;
		correct = 32'b00001011010001100010000110110000;
		#400 //-3.5692643e-24 * -93537224.0 = 3.8158757e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011010101110000010001000111;
		b = 32'b10010110000010101100101011000001;
		correct = 32'b01110100110001100100110000110111;
		#400 //-14091335.0 * -1.1211529e-25 = 1.2568611e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100010101011011010000101010101;
		b = 32'b11011000111000101010001000110110;
		correct = 32'b10001001010001000010000011101010;
		#400 //4.706256e-18 * -1993490500000000.0 = -2.3608118e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101100110101110010001010000111;
		b = 32'b10001001101010111110100010101001;
		correct = 32'b01100010101000000010111101101110;
		#400 //-6.114501e-12 * -4.1385545e-33 = 1.4774484e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010101001110110001110001111001;
		b = 32'b11111011101100001110011001100011;
		correct = 32'b10011001000001110110001101111011;
		#400 //12858185000000.0 * -1.8370341e+36 = -6.999426e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001011001001110110011110111011;
		b = 32'b10001111111111011110010100111001;
		correct = 32'b10111010101010001100101011111001;
		#400 //3.2241068e-32 * -2.503602e-29 = -0.0012877873
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110100001011100010011001110011;
		b = 32'b10110100101001101111111110000001;
		correct = 32'b11111111000001010111101101100000;
		#400 //5.51904e+31 * -3.1105813e-07 = -1.7742792e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011000010111000110000101101111;
		b = 32'b00110100001010111001001010000000;
		correct = 32'b11100011101001000110100110111101;
		#400 //-969244100000000.0 * 1.5978912e-07 = -6.0657705e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000110011000101111001001000011;
		b = 32'b00110101100100000110000101010101;
		correct = 32'b01010000010010010011001011101000;
		#400 //14524.565 * 1.0757163e-06 = 13502226000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011110011001110100100101001111;
		b = 32'b00111110010000110010100001101011;
		correct = 32'b01011111100101111011001000101000;
		#400 //4.1664847e+18 * 0.19058387 = 2.1861686e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011101001011100000110101111100;
		b = 32'b11001111011011010010001011111011;
		correct = 32'b00001101001110111110010111011111;
		#400 //-2.303568e-21 * -3978492700.0 = 5.790052e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110100001110000010010011001011;
		b = 32'b10111110011010100010010011001011;
		correct = 32'b11110101010010010101010100101101;
		#400 //5.8357475e+31 * -0.22865598 = -2.5521954e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001101111110100111001010000101;
		b = 32'b10000111011011110000100000001000;
		correct = 32'b11000110000001100001110011111010;
		#400 //1.5435009e-30 * -1.7982722e-34 = -8583.244
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010110111000010001000110110001;
		b = 32'b00110100100010011000110011011010;
		correct = 32'b01100001110100010111000101000010;
		#400 //123733050000000.0 * 2.5620722e-07 = 4.8294132e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110000010001010101100000100011;
		b = 32'b11010100100101011010100111110111;
		correct = 32'b01011011001010001100011101010011;
		#400 //-2.443004e+29 * -5142413300000.0 = 4.7506955e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000001001010100011101101111100;
		b = 32'b00100101011111000001001100101101;
		correct = 32'b10011011001011001110001000010001;
		#400 //-3.1266747e-38 * 2.1864013e-16 = -1.4300553e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111001100001111100000000100100;
		b = 32'b11110100110111000011100010111000;
		correct = 32'b00000100000111011100111000101100;
		#400 //-0.00025892362 * -1.39581995e+32 = 1.854993e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011110010001011001110101011011;
		b = 32'b01000010110010001110100101111101;
		correct = 32'b01011010111110111100110001101010;
		#400 //3.5599094e+18 * 100.45603 = 3.5437487e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110110101001010110010010001001;
		b = 32'b00111001100110000110010111000010;
		correct = 32'b01111100100010101110101000110001;
		#400 //1.6772814e+33 * 0.00029067515 = 5.7702955e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011010100001000010100001110100;
		b = 32'b10101001111010001010100100010001;
		correct = 32'b00110000000100010110101001100101;
		#400 //-5.4659276e-23 * -1.0332198e-13 = 5.290189e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010001000110111000000101100101;
		b = 32'b01001101000001010000010000001001;
		correct = 32'b11000011100101011010010001000011;
		#400 //-41743176000.0 * 139477140.0 = -299.2833
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110000011111100111001101011100;
		b = 32'b10001111111010110011000011111000;
		correct = 32'b11100000000010100111101101001110;
		#400 //9.25686e-10 * -2.3191651e-29 = -3.991462e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100010001000010101101111100110;
		b = 32'b10111101100010000101010111010100;
		correct = 32'b00100100000101110111111001101010;
		#400 //-2.186822e-18 * -0.066569954 = 3.2849982e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111110111111000100001110011101;
		b = 32'b00101001011111100010101101010100;
		correct = 32'b11010100111111100001010011000110;
		#400 //-0.49270335 * 5.643691e-14 = -8730161700000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111011110101110000111111100110;
		b = 32'b01100011111011101010100110001111;
		correct = 32'b01010111011001101010111101110001;
		#400 //2.2333326e+36 * 8.805086e+21 = 253641190000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001101101110101100110110011101;
		b = 32'b11000000100100001110010100010101;
		correct = 32'b00001100101001010000010110010100;
		#400 //-1.1512635e-30 * -4.527964 = 2.5425632e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111100111101101001101001001010;
		b = 32'b00110101011111000111011011110011;
		correct = 32'b01000110111110100000111001010011;
		#400 //0.030102868 * 9.405041e-07 = 32007.162
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001110000100100100001110101001;
		b = 32'b01000111111100111000001101110001;
		correct = 32'b11000101100110011100001110100101;
		#400 //-613476900.0 * 124678.88 = -4920.4556
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010101100000111010111001110010;
		b = 32'b00111000110011000111111100110110;
		correct = 32'b00011100001001001101100010000010;
		#400 //5.3185705e-26 * 9.751173e-05 = 5.454288e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110111000010000111100101110010;
		b = 32'b10111010001010011011011111010011;
		correct = 32'b10111100010011011101101100010101;
		#400 //8.134508e-06 * -0.00064742303 = -0.01256444
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110111001101100110101001101100;
		b = 32'b11001000010101110010000011101101;
		correct = 32'b01101110010110010001001001110110;
		#400 //-3.6998302e+33 * -220291.7 = 1.6795141e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110110101001110011111111101010;
		b = 32'b01011100000001101110110111110010;
		correct = 32'b00011010000111101010100100001100;
		#400 //4.9844284e-06 * 1.5191708e+17 = 3.281019e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100101010110110000100001111100;
		b = 32'b00010011011110001111011011100110;
		correct = 32'b01010001011000010011100100001101;
		#400 //1.8998097e-16 * 3.1423731e-27 = 60457800000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010101101011100001111110111111;
		b = 32'b10101100110010011001100111010110;
		correct = 32'b10101000010111010001101111011101;
		#400 //7.0328127e-26 * -5.729843e-12 = -1.2274006e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010101110110001100000101110111;
		b = 32'b11001101111100000011011000111010;
		correct = 32'b10000111011001110000000010010010;
		#400 //8.754694e-26 * -503760700.0 = -1.7378676e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000110010001101110100010011110;
		b = 32'b10111011011110111100110010001110;
		correct = 32'b01001010010010100011101000101010;
		#400 //-12730.154 * -0.0038421485 = 3313290.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101000111000010100011001001000;
		b = 32'b10001101100100010011110001100101;
		correct = 32'b11011010110001101000101000111110;
		#400 //2.5010498e-14 * -8.950854e-31 = -2.7942022e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111111101110000100000110111100;
		b = 32'b11101001011101100111111000011101;
		correct = 32'b10010101101111110101110100011001;
		#400 //1.439506 * -1.8624457e+25 = -7.729117e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000100000011010000001011100111;
		b = 32'b10000001011001010000001000010011;
		correct = 32'b01000010000111011010000110101101;
		#400 //-1.6575803e-36 * -4.2062145e-38 = 39.407887
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101001010100010100100100010111;
		b = 32'b01011010111111000100100001101011;
		correct = 32'b11001101110101000101111001111110;
		#400 //-1.5813166e+25 * 3.550566e+16 = -445370300.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011011001101111111000000001011;
		b = 32'b01100000101011100111101010011100;
		correct = 32'b00111010000001101111000001100101;
		#400 //5.177385e+16 * 1.0058026e+20 = 0.0005147516
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001110000111101001111101010110;
		b = 32'b01010111111100011000011011110001;
		correct = 32'b10110101101010000010000010100000;
		#400 //-665310600.0 * 531123740000000.0 = -1.252647e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100001110001111101110011011101;
		b = 32'b10111110011110011000100001101111;
		correct = 32'b00100010110011010000101011100011;
		#400 //-1.3543227e-18 * -0.24368452 = 5.557689e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011100010110101101010001000101;
		b = 32'b10011100111100100111101011001001;
		correct = 32'b10111110111001110000011111100100;
		#400 //7.24045e-22 * -1.6045956e-21 = -0.45123208
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100000111101010101001111111001;
		b = 32'b01100100000010011010011010001100;
		correct = 32'b00111100011001000010000011010110;
		#400 //1.4142197e+20 * 1.015682e+22 = 0.013923844
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011101111011001110100111000000;
		b = 32'b10101011000011111101110010101000;
		correct = 32'b10110010010100101100101010100000;
		#400 //6.271037e-21 * -5.111003e-13 = -1.226968e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001001000000000111101110101101;
		b = 32'b00001101000100111010111101010010;
		correct = 32'b10111011010111101011011100011110;
		#400 //-1.5465592e-33 * 4.5508906e-31 = -0.0033983658
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111000010111011000110010001011;
		b = 32'b10000100010110110011010110010010;
		correct = 32'b01110011100000010101110111000000;
		#400 //-5.2821397e-05 * -2.5767925e-36 = 2.0498894e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100100111010000101010011100010;
		b = 32'b01001111010111001010100000000001;
		correct = 32'b00010101000001101100010111010000;
		#400 //1.0075776e-16 * 3701997800.0 = 2.721713e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100100110010111011010001000001;
		b = 32'b01000010010100110110111001001011;
		correct = 32'b00100001111101101010010011111111;
		#400 //8.834258e-17 * 52.857708 = 1.6713283e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000001101001111011110001100010;
		b = 32'b10111010001001100010001011111101;
		correct = 32'b11000111000000010011101101101011;
		#400 //20.966984 * -0.0006337611 = -33083.418
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100011100100011000101111110100;
		b = 32'b00110011010010011111010000001100;
		correct = 32'b11101111101110000111111101110100;
		#400 //-5.369725e+21 * 4.702092e-08 = -1.1419865e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001000011000000010000101100111;
		b = 32'b11010101110011000110001010011011;
		correct = 32'b10110010000011000101110110101001;
		#400 //229509.61 * -28090485000000.0 = -8.170368e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111010000010000110010011011010;
		b = 32'b01100001000100001001011101101101;
		correct = 32'b11011000011100010111110001110111;
		#400 //-1.7704947e+35 * 1.6670266e+20 = -1062067500000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010010001001110000010100111101;
		b = 32'b11100111000110010010011100101110;
		correct = 32'b10101010100010111001011100000100;
		#400 //179336860000.0 * -7.232448e+23 = -2.4796148e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101110010111010011000010110101;
		b = 32'b11001010001010111101010010011011;
		correct = 32'b10100011101001001100010011100011;
		#400 //5.0292843e-11 * -2815270.8 = -1.78643e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010000110011101100011001010100;
		b = 32'b10010001100101101111001110101100;
		correct = 32'b11111110101011110101010111001100;
		#400 //27752833000.0 * -2.3816002e-28 = -1.1653019e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010110010111011010000101011011;
		b = 32'b11001000010111110000100011011001;
		correct = 32'b10001101011111100110001101100000;
		#400 //1.7903153e-25 * -228387.39 = -7.838941e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011110010100110010111111010110;
		b = 32'b10111100010010101101110010000011;
		correct = 32'b11100001100001010100000011001111;
		#400 //3.8044042e+18 * -0.012381676 = -3.0726086e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000110101000100100000110010000;
		b = 32'b00101000101110101011010001000101;
		correct = 32'b10011101010111100111101001011011;
		#400 //-6.103396e-35 * 2.0728328e-14 = -2.9444712e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110110100011101010100101111011;
		b = 32'b11010111101110010000011010100111;
		correct = 32'b10011110010001010110001010111100;
		#400 //4.25166e-06 * -406876450000000.0 = -1.0449511e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010101101001110111001001000101;
		b = 32'b00111101001010101100111001111110;
		correct = 32'b10010111111110101111011010111001;
		#400 //-6.763105e-26 * 0.041700833 = -1.6218153e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111101100110001100000101100100;
		b = 32'b10000011010011100000001011111111;
		correct = 32'b11111001101111011101001000111011;
		#400 //0.07458761 * -6.05414e-37 = -1.2320101e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001010101100011010111101001110;
		b = 32'b10111100111000001100101011011110;
		correct = 32'b10001101010010100101101000111011;
		#400 //1.7110422e-32 * -0.027440485 = -6.2354667e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101010001101101110111100101110;
		b = 32'b00001101011101010011010000100000;
		correct = 32'b11011100001111101111110100101100;
		#400 //-1.624783e-13 * 7.5559197e-31 = -2.1503444e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010111100101010000000111100110;
		b = 32'b10111100111001101001100001110110;
		correct = 32'b01011010001001010110110001100011;
		#400 //-327670770000000.0 * -0.02814887 = 1.1640636e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011101011101011100000011110010;
		b = 32'b10001100110011010010011101010111;
		correct = 32'b11010000000110010101010011001110;
		#400 //3.252523e-21 * -3.1608928e-31 = -10289887000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111000111100101001111011110100;
		b = 32'b10111110101001010011011001110001;
		correct = 32'b10111001101110111111100100000101;
		#400 //0.000115690666 * -0.32268098 = -0.00035852953
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000100010101001000011011011110;
		b = 32'b00101000110100111100000100100100;
		correct = 32'b11011011000000000111011110000101;
		#400 //-850.1073 * 2.3509467e-14 = -3.616021e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100011111100011011010100100;
		b = 32'b01010000010011100110100011000100;
		correct = 32'b00110011100111011010010100001010;
		#400 //1016.85376 * 13851890000.0 = 7.3409026e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111100000111010010101101001;
		b = 32'b00100000100010101001111010100101;
		correct = 32'b01100110011100110001111100010001;
		#400 //67402.82 * 2.3483091e-19 = 2.8702703e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110100010101010011000011101100;
		b = 32'b10101110001011111001000011101101;
		correct = 32'b01000101100110110110111001100110;
		#400 //-1.9854969e-07 * -3.9919113e-11 = 4973.8
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100100101101010111111000001001;
		b = 32'b11111100000000011011011110110001;
		correct = 32'b10101000001100110001011011011001;
		#400 //2.678354e+22 * -2.694128e+36 = -9.94145e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100100111100010101011111111000;
		b = 32'b11100110001111110011110100110101;
		correct = 32'b10111110001000011000100100110011;
		#400 //3.5616033e+22 * -2.2577527e+23 = -0.15774994
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101101010111001010011011000110;
		b = 32'b01010011011001101000100010001000;
		correct = 32'b01011001011101010000011011001001;
		#400 //4.26802e+27 * 990133100000.0 = 4310551900000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011111000111010001001011100;
		b = 32'b10111011011001011101110011010100;
		correct = 32'b01001111111111011000010010101010;
		#400 //-29836472.0 * -0.003507425 = 8506660000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011110100101101010100011000001;
		b = 32'b11000100010100010100101011010101;
		correct = 32'b00011001101110000100100000100001;
		#400 //-1.5951663e-20 * -837.16925 = 1.9054287e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011111000100010011111010100100;
		b = 32'b10101100110110110100001111101011;
		correct = 32'b11110001101010011001010000001100;
		#400 //1.0465983e+19 * -6.2318948e-12 = -1.6794222e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100101010001010101010101011010;
		b = 32'b01011010111101010000110110001101;
		correct = 32'b11001001110011100010011000010011;
		#400 //-5.824254e+22 * 3.4488134e+16 = -1688770.4
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101110011000111110001000100011;
		b = 32'b11010111010001001011110111010010;
		correct = 32'b01010110100101000100001011001010;
		#400 //-1.763162e+28 * -216319550000000.0 = 81507290000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111011111010010010110101010001;
		b = 32'b00101000111111110100001011101010;
		correct = 32'b01010010011010011101101000001011;
		#400 //0.007115998 * 2.8339706e-14 = 251096380000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100011000011011100011111101110;
		b = 32'b00001010110010001011111101001000;
		correct = 32'b01010111101101001100110111011110;
		#400 //7.685962e-18 * 1.9331251e-32 = 397592570000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001110011000000110110100000100;
		b = 32'b10010011101100000000001001101010;
		correct = 32'b11111010001000110011010111000110;
		#400 //941310200.0 * -4.4431027e-27 = -2.1185876e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111011110010010110101001001100;
		b = 32'b11101000010011011100010011011101;
		correct = 32'b11010010111110101001010101011010;
		#400 //2.0916153e+36 * -3.8868665e+24 = -538123760000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010011011000111010110010111001;
		b = 32'b10101001000010001010111110110011;
		correct = 32'b10101001110101010011010011000100;
		#400 //2.8736587e-27 * -3.035046e-14 = -9.4682535e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100010000101111110101100000110;
		b = 32'b11011111001001010101001101011101;
		correct = 32'b11000010011010110011110100101001;
		#400 //7.005984e+20 * -1.1912968e+19 = -58.809727
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100100110011110000101101001010;
		b = 32'b10010001001010101000011010011000;
		correct = 32'b11010011000110110110100101010001;
		#400 //8.9791064e-17 * -1.345211e-28 = -667486850000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110101111100010111100100010000;
		b = 32'b11000010000001010011101000011110;
		correct = 32'b11110011011001111111111110111100;
		#400 //6.1220653e+32 * -33.306755 = -1.8380851e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110110011101001001100000111011;
		b = 32'b00001100011011110000100011101101;
		correct = 32'b01101001100000101111101000101001;
		#400 //3.6447443e-06 * 1.8414576e-31 = 1.9792713e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100110001001110001000010011011;
		b = 32'b10110101000110110010100000011001;
		correct = 32'b11110000100010011101001011110000;
		#400 //1.9723538e+23 * -5.780035e-07 = -3.4123563e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010011100100010110101000110100;
		b = 32'b00100000100000100010011100011010;
		correct = 32'b11110010100011110000001001111010;
		#400 //-1249104100000.0 * 2.2048732e-19 = -5.665197e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101011110010010101110110100010;
		b = 32'b10111010100110111010110010001011;
		correct = 32'b01110000101001011001000110110110;
		#400 //-4.868725e+26 * -0.0011876983 = 4.0992944e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101110010001100011100001110111;
		b = 32'b01010001101010101100100001100110;
		correct = 32'b10011100000101001001000001111000;
		#400 //-4.507014e-11 * 91688320000.0 = -4.9155814e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011011011101011100111110000110;
		b = 32'b01101110011111101111011100001101;
		correct = 32'b10101100011101101100111011110110;
		#400 //-6.9189544e+16 * 1.9726965e+28 = -3.507359e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000010110001011010110001110100;
		b = 32'b00111011001011110010101011100001;
		correct = 32'b11000111000100000111001000100110;
		#400 //-98.83682 * 0.0026728439 = -36978.15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100101001110111110110110001101;
		b = 32'b10111110000110101111110001110100;
		correct = 32'b01100110100110110011010010111011;
		#400 //-5.5466536e+22 * -0.15135366 = 3.6646976e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100000110010010001001100011110;
		b = 32'b00101001010000100111001111100101;
		correct = 32'b01110111000001000101101111100101;
		#400 //1.1591166e+20 * 4.3177176e-14 = 2.6845587e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000010100011110110111001111001;
		b = 32'b00000000101111101100100011000011;
		correct = 32'b11000001010000000111010111110011;
		#400 //-2.107537e-37 * 1.7520764e-38 = -12.028796
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010110110001001111001111010111;
		b = 32'b11000001101100111110000011010001;
		correct = 32'b11010100100011000010011001100011;
		#400 //108275780000000.0 * -22.484774 = -4815515500000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101011001100011110100010001001;
		b = 32'b10111101101100011000010011010101;
		correct = 32'b11101101000000000100011111100100;
		#400 //2.1507799e+26 * -0.08667914 = -2.481312e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001101101000100010010100101001;
		b = 32'b00011000011111110010101000011110;
		correct = 32'b01110100101000101010110100010011;
		#400 //340043040.0 * 3.2979241e-24 = 1.0310821e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101111110011101100010000111111;
		b = 32'b01010111011111001000001001101011;
		correct = 32'b00010111110100011001111111110100;
		#400 //3.7610623e-10 * 277637070000000.0 = 1.3546686e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100000001100100001000001101010;
		b = 32'b10011011110101111000100100111011;
		correct = 32'b11000011110100110111111001000011;
		#400 //1.5082617e-19 * -3.565745e-22 = -422.98642
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111100011001001100011111110011;
		b = 32'b01010010101001111100101100111110;
		correct = 32'b01101001001011101000011000000001;
		#400 //4.7515965e+36 * 360334700000.0 = 1.3186619e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001100010101100000010100010010;
		b = 32'b10111010100111110101110110010101;
		correct = 32'b11010001001010111110010111000000;
		#400 //56104010.0 * -0.0012158627 = -46143373000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011001100010000000010110111001;
		b = 32'b10011001011111101011111111000100;
		correct = 32'b10111111100010001011000010110110;
		#400 //1.4064382e-23 * -1.3170219e-23 = -1.0678928
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111111110100100111010011111111;
		b = 32'b11110001110000011111000100101110;
		correct = 32'b00001101100010101110011001010010;
		#400 //-1.6441954 * -1.9207096e+30 = 8.560354e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000011101101000001010100010001;
		b = 32'b00101000001100010100100101111010;
		correct = 32'b11011011000000100000010010100111;
		#400 //-360.16458 * 9.8414065e-15 = -3.6596862e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001011010000111011011101001000;
		b = 32'b10101110111101100101111000001000;
		correct = 32'b00011011110010110101111001000100;
		#400 //-3.769352e-32 * -1.1203488e-10 = 3.364445e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111000100000100011101111111111;
		b = 32'b00111100010000101000010110010011;
		correct = 32'b01111011101010110110010100001001;
		#400 //2.1131733e+34 * 0.011872667 = 1.779864e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001000101011010001011011101100;
		b = 32'b10110001010110111111011101011001;
		correct = 32'b10010110110010010111000110111001;
		#400 //1.0417448e-33 * -3.2009295e-09 = -3.254507e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100101111110011110101000101101;
		b = 32'b00010001111011111100011110101001;
		correct = 32'b01010011100001010110100100000011;
		#400 //4.3353298e-16 * 3.7830601e-28 = 1145984900000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000001011110000110111100111011;
		b = 32'b00001100110011000000100110111110;
		correct = 32'b00110100000110111101100111110101;
		#400 //4.563021e-38 * 3.143704e-31 = 1.4514792e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011110010011100011000010010110;
		b = 32'b10010011010110101001011001011011;
		correct = 32'b11001010011100010111101100000101;
		#400 //1.09155965e-20 * -2.75896e-27 = -3956417.2
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010010001001110110111011010010;
		b = 32'b10111011101110100110111100011011;
		correct = 32'b11010101111001011110100010101000;
		#400 //179779700000.0 * -0.0056895143 = -31598427000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000011110001100001101110110111;
		b = 32'b11001000001110100000100110000000;
		correct = 32'b00111011000010000100111000101101;
		#400 //-396.21652 * -190502.0 = 0.002079855
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001110011100111101110000001100;
		b = 32'b10111111010101010001101000101100;
		correct = 32'b00001110100100100111100101110011;
		#400 //-3.0058011e-30 * -0.8324306 = 3.610873e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111110110010010101111100110110;
		b = 32'b11000001001111101111100000110110;
		correct = 32'b01111101000001101111100011101010;
		#400 //-1.338346e+38 * -11.935598 = 1.1213062e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101101001010010001000101010100;
		b = 32'b10111111100011001111010001001010;
		correct = 32'b10101101000110011000011110011010;
		#400 //9.610385e-12 * -1.1012051 = -8.727153e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111000001110001000010001001010;
		b = 32'b00100100110101000001101010110011;
		correct = 32'b11010010110111101011010000000000;
		#400 //-4.3992222e-05 * 9.1985574e-17 = -478251320000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010111010101000111101101110110;
		b = 32'b10111101000000111110101001111000;
		correct = 32'b01011001110011100010110010111110;
		#400 //-233626730000000.0 * -0.03220603 = 7254130000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101010100100101101010001110000;
		b = 32'b00101110100011100011011001011111;
		correct = 32'b01111011100001000010011111101111;
		#400 //8.875319e+25 * 6.4670706e-11 = 1.3723863e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101101000001100010100000000011;
		b = 32'b01010001110111111010001110101101;
		correct = 32'b00011010100110011001000110011000;
		#400 //7.6259025e-12 * 120065470000.0 = 6.3514536e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010000000110000101110000001101;
		b = 32'b00101010011110011011011010000011;
		correct = 32'b01100101000111000011001000010000;
		#400 //10224678000.0 * 2.2178964e-13 = 4.610079e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111011110000011011101100110100;
		b = 32'b00110011011111110101011111101011;
		correct = 32'b11000111110000100011101010111010;
		#400 //-0.005912209 * 5.9451775e-08 = -99445.45
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001100110111110110100001010111;
		b = 32'b10001000011100110011111000101011;
		correct = 32'b01000011111010110001111111011100;
		#400 //-3.4421387e-31 * -7.319823e-34 = 470.2489
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101111010100011111010100000100;
		b = 32'b10001111001010011100010011001011;
		correct = 32'b11011111100111100100110011111011;
		#400 //1.9095486e-10 * -8.370244e-30 = -2.2813536e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101101001111011110000000110100;
		b = 32'b00111011110101111010101100001011;
		correct = 32'b10110000111000010110001001011111;
		#400 //-1.0793189e-11 * 0.006581669 = -1.6398863e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101110111111010101011111010111;
		b = 32'b10110000001100110011101100110101;
		correct = 32'b11111110001101001110110110000100;
		#400 //3.920295e+28 * -6.520396e-10 = -6.0123573e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000001010100010111100011011001;
		b = 32'b00111111011011011111010001011010;
		correct = 32'b00000001011000010101101110001010;
		#400 //3.847394e-38 * 0.92950976 = 4.139165e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100111101100000001000110100110;
		b = 32'b01111100111110100100110101101100;
		correct = 32'b10101010001101000001001110100110;
		#400 //-1.6629241e+24 * 1.0397156e+37 = -1.5994028e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111110011010111110010100100000;
		b = 32'b11110101010101000111011000001000;
		correct = 32'b11001000100011100001111000111100;
		#400 //7.8389566e+37 * -2.6932639e+32 = -291057.88
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011010101100010110011010010111;
		b = 32'b00100010001000100001101001101100;
		correct = 32'b11111000000011000001010001001001;
		#400 //-2.4966935e+16 * 2.1969082e-18 = -1.1364578e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110110101100110010000011011111;
		b = 32'b01101111101100100101110001101100;
		correct = 32'b01000110100000001000110011111011;
		#400 //1.8165778e+33 * 1.1040013e+29 = 16454.49
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111111110011010010011111110011;
		b = 32'b10001010101110110111100011011001;
		correct = 32'b01110100100011000001001011110110;
		#400 //-1.6027817 * -1.8052903e-32 = 8.878249e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101010100110001101011111111110;
		b = 32'b00000001000000100001001100100110;
		correct = 32'b01101001000101100110011111011110;
		#400 //2.71505e-13 * 2.3890967e-38 = 1.1364336e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011110101101100011101000111001;
		b = 32'b11001000000110100000001110011110;
		correct = 32'b01010110000101110111001010100111;
		#400 //-6.565435e+18 * -157710.47 = 41629670000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100110011011100001100001010101;
		b = 32'b11100000011101011101101110101110;
		correct = 32'b11000101011101111110101010101100;
		#400 //2.8109302e+23 * -7.086378e+19 = -3966.667
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100110010010101011100001010001;
		b = 32'b00100000111111111111100101000011;
		correct = 32'b01000100110010101011110110100111;
		#400 //7.0332624e-16 * 4.3363628e-19 = 1621.9266
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100011010000000001000011011010;
		b = 32'b10010110101110010110010001110110;
		correct = 32'b01001100000001001001101110000101;
		#400 //-1.0411909e-17 * -2.9951762e-25 = 34762260.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100011001011110000000101001111;
		b = 32'b00111011000010101010100110100000;
		correct = 32'b11100111101000011000110001000101;
		#400 //-3.2282745e+21 * 0.0021158233 = -1.525777e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110100111111110101000000001000;
		b = 32'b10101101000011110110001101001011;
		correct = 32'b01000111011000111110100111010101;
		#400 //-4.7555682e-07 * -8.150656e-12 = 58345.832
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011001101011110011111100110111;
		b = 32'b11000001100010100011100111101100;
		correct = 32'b01010111101000100100100000100101;
		#400 //-6165953300000000.0 * -17.278282 = 356861500000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001000100101010011100100100010;
		b = 32'b00111101000101100111010100101001;
		correct = 32'b10001010111111011110011001001010;
		#400 //-8.981043e-34 * 0.036732826 = -2.4449639e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101010001110111111010111000100;
		b = 32'b01001111011110011010001000011010;
		correct = 32'b10011010010000001100000011111101;
		#400 //-1.6694204e-13 * 4188150300.0 = -3.9860564e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010111101001100110011000011101;
		b = 32'b11111100011111111001111110100111;
		correct = 32'b00011010101001101010010011010101;
		#400 //-365915000000000.0 * -5.3090953e+36 = 6.892229e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001010001001101101111011111101;
		b = 32'b10110111101101110001010111011010;
		correct = 32'b10010001111010010101010000001001;
		#400 //8.034549e-33 * -2.1825475e-05 = -3.681271e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010001000111000000101000011011;
		b = 32'b11011101010101100101000011010100;
		correct = 32'b10110011001110100110001110011001;
		#400 //41886527000.0 * -9.6519226e+17 = -4.3397083e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011100001011011011000111000110;
		b = 32'b11011011010101000001001011111001;
		correct = 32'b01000000010100011010101111000001;
		#400 //-1.9556254e+17 * -5.9693556e+16 = 3.276108
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101011101011010000110101110011;
		b = 32'b00111110001111010001011000111000;
		correct = 32'b11101100111010100100101010100111;
		#400 //-4.1841536e+26 * 0.18465507 = -2.2659294e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111100011110111111001111010111;
		b = 32'b11101111000111000101110110001110;
		correct = 32'b00001100110011100011111101000010;
		#400 //-0.01537796 * -4.839276e+28 = 3.1777397e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100110010100101011011001010100;
		b = 32'b10101111110101110010000011110100;
		correct = 32'b10110101111110101011111010010011;
		#400 //7.3105487e-16 * -3.9131687e-10 = -1.8681916e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011111100011010000111001100011;
		b = 32'b00101100011000000100010010001010;
		correct = 32'b11110010101000010000001110111111;
		#400 //-2.032834e+19 * 3.1870361e-12 = -6.378447e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100100011110111101010011000011;
		b = 32'b01001100110101011000100101011011;
		correct = 32'b00010111000101101111010001110010;
		#400 //5.4607165e-17 * 111954650.0 = 4.8776147e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110100110101110110000010101;
		b = 32'b11010111011100111010101011100011;
		correct = 32'b10100110101000101100001101011011;
		#400 //0.3025824 * -267915280000000.0 = -1.1293959e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101101110111100000000111101001;
		b = 32'b00011010001100010010100100000010;
		correct = 32'b11010011001000000110011100010001;
		#400 //-2.5239326e-11 * 3.6635868e-23 = -688923930000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010000101011101011001111011011;
		b = 32'b11000100100000100101000010100000;
		correct = 32'b01001011101010111001100101011111;
		#400 //-23448180000.0 * -1042.5195 = 22491838.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110011110100101111010010111111;
		b = 32'b01000001000001101110010100000100;
		correct = 32'b01110010010010000010110010000011;
		#400 //3.3427319e+31 * 8.430912 = 3.964852e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010001101001100000011100101000;
		b = 32'b10111011010100001011101100010111;
		correct = 32'b10010101110010111010000001101100;
		#400 //2.6194592e-28 * -0.0031849795 = -8.224415e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100000101000101000011101101001;
		b = 32'b10010001010101010110110101100000;
		correct = 32'b11001110110000101111001011101100;
		#400 //2.7533474e-19 * -1.6836441e-28 = -1635350000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110100101001010000101101100110;
		b = 32'b00010100011010001101000110101100;
		correct = 32'b01011111101101010111101000111001;
		#400 //3.0741938e-07 * 1.1754357e-26 = 2.6153654e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101101011010000110000101010001;
		b = 32'b00000010101111011001110100101011;
		correct = 32'b11101010000111001101111010011101;
		#400 //-1.3209282e-11 * 2.7861264e-37 = -4.7410922e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110011000111100001010100101101;
		b = 32'b10111110000111101001100010111010;
		correct = 32'b01110100011111110010101110101000;
		#400 //-1.2524603e+31 * -0.15487948 = 8.086677e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011001110110000100011010101010;
		b = 32'b10100001001010001110110100011110;
		correct = 32'b11111000001000111110000011010011;
		#400 //7609536400000000.0 * -5.7234436e-19 = -1.3295381e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101011101100010010000101001000;
		b = 32'b10100110111001110001011101110000;
		correct = 32'b01000100010001000011100011011111;
		#400 //-1.2585844e-12 * -1.6035198e-15 = 784.8886
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011111001000111010010011000110;
		b = 32'b11011011011101011010010010010110;
		correct = 32'b00000011001010101000101100011011;
		#400 //-3.465289e-20 * -6.9142333e+16 = 5.0118195e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001001010111101001001011101011;
		b = 32'b10100101110110000000111110101100;
		correct = 32'b10100011000000111101101110111000;
		#400 //2.6791358e-33 * -3.7480647e-16 = -7.1480515e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000101101111011010010110000100;
		b = 32'b10011000000001110111100011000101;
		correct = 32'b10101101001100110010111111010110;
		#400 //1.7834275e-35 * -1.7509314e-24 = -1.0185594e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100100101110110011100000010001;
		b = 32'b00100111001001001111101100011110;
		correct = 32'b01111101000100010100000011011100;
		#400 //2.762865e+22 * 2.2895703e-15 = 1.2067177e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010011100001110011000011100;
		b = 32'b00111101011010101010100011111110;
		correct = 32'b10111100100000110110011100101110;
		#400 //-0.00091895624 * 0.05729007 = -0.01604041
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111010011101101000111001111111;
		b = 32'b11010011101111101001011001110011;
		correct = 32'b01100110001001011001011011010001;
		#400 //-3.200488e+35 * -1637135800000.0 = 1.9549314e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111100101010010010101010000010;
		b = 32'b01100001010110101110101000000110;
		correct = 32'b10011010110001011101001011111100;
		#400 //-0.020650152 * 2.5239084e+20 = -8.1818154e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011010001101001010000000111110;
		b = 32'b00011011000010101111000000010110;
		correct = 32'b00111110101001100110011111111111;
		#400 //3.735257e-23 * 1.1492668e-22 = 0.32501218
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000110101111000010110000110;
		b = 32'b10100000110100100101011010110101;
		correct = 32'b01001111100000110010011101101101;
		#400 //-1.5681259e-09 * -3.5632762e-19 = 4400798000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000010101111101100111010000010;
		b = 32'b11101101111111110100101010000110;
		correct = 32'b10010100001111110101011000100101;
		#400 //95.403336 * -9.8760964e+27 = -9.660025e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011100011110111100101001001000;
		b = 32'b00001010001001100010111011000000;
		correct = 32'b11010001110000011111000000100111;
		#400 //-8.3310376e-22 * 8.001402e-33 = -104119720000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011100111011100010100101111000;
		b = 32'b01100000100100010110000010010010;
		correct = 32'b00111011110100011011000110101011;
		#400 //5.3629312e+17 * 8.380427e+19 = 0.0063993535
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001101000011100100011001000011;
		b = 32'b10111001010101110010000000111101;
		correct = 32'b00010011001010010100111010000100;
		#400 //-4.3841703e-31 * -0.00020516007 = 2.136951e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111001001011010111100000100000;
		b = 32'b10111110000110011100100001101010;
		correct = 32'b10111010100100000110001011000100;
		#400 //0.00016543316 * -0.15017858 = -0.0011015763
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111101010100110000001010111111;
		b = 32'b11010110010100010010000010001000;
		correct = 32'b10100110100000010010011100100110;
		#400 //0.05151629 * -57484413000000.0 = -8.961784e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100110111010110000101001011000;
		b = 32'b10110111010101001001101011000010;
		correct = 32'b01101111000011011000000111110111;
		#400 //-5.5497347e+23 * -1.2672217e-05 = 4.3794504e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100111001111010010010010010010;
		b = 32'b01100101001101100001100010011111;
		correct = 32'b10000001100001001111010000001011;
		#400 //-2.6248844e-15 * 5.3745305e+22 = -4.8839326e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010011001010100001110111100010;
		b = 32'b10001101101010011100010010100101;
		correct = 32'b01000101000000000100001101001000;
		#400 //-2.147175e-27 * -1.046277e-30 = 2052.205
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110001000001010100101111001010;
		b = 32'b11101111000101111111000101101010;
		correct = 32'b00000001011000001001010100110010;
		#400 //-1.9397128e-09 * -4.702409e+28 = 4.1249345e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110111101001010010000101100110;
		b = 32'b01110001110100011101010000011101;
		correct = 32'b11000101010010010111011101100100;
		#400 //-6.6984874e+33 * 2.0780415e+30 = -3223.462
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111100101000101010010000011110;
		b = 32'b01000110100100011111010100101111;
		correct = 32'b00110101100011101010000101110111;
		#400 //0.019853648 * 18682.592 = 1.0626817e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000011001110010000101010110000;
		b = 32'b10111001011001100010101110000001;
		correct = 32'b11001001010011011100111010110101;
		#400 //185.04175 * -0.00021950716 = -842987.3
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111001001000101110111000110111;
		b = 32'b10100100011001110110101111110101;
		correct = 32'b11010100001101000011110000010011;
		#400 //0.00015538266 * -5.0181584e-17 = -3096408000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110011000011001111111001011101;
		b = 32'b01110110011110100001010110011010;
		correct = 32'b10111100000100000101010000101000;
		#400 //-1.1170664e+31 * 1.2680785e+33 = -0.008809127
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101100111011000111100010100010;
		b = 32'b01001111000000001111001001101010;
		correct = 32'b01011101011010101011110000010100;
		#400 //2.2870093e+27 * 2163370500.0 = 1.057151e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001100010111000110111101101000;
		b = 32'b10010011000101111111110110001101;
		correct = 32'b11111000101110011010010000101101;
		#400 //57785760.0 * -1.918389e-27 = -3.0122025e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100010110101110001001110111101;
		b = 32'b00101100010011011100010010011001;
		correct = 32'b11110110000001011100101001110101;
		#400 //-1.9837361e+21 * 2.9241386e-12 = -6.784002e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101011011110101110011000000100;
		b = 32'b11011111010001010000101111011010;
		correct = 32'b00001011101000101111101101100111;
		#400 //-8.9137053e-13 * -1.4198682e+19 = 6.27784e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101101010001101111001101100011;
		b = 32'b11011011000101110100000000110010;
		correct = 32'b11010001101010000101111000001100;
		#400 //3.8482668e+27 * -4.2573305e+16 = -90391540000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101001110101011010101001010110;
		b = 32'b11100000101010000000101110000100;
		correct = 32'b00001000101000101011111111000100;
		#400 //-9.488649e-14 * -9.687134e+19 = 9.795104e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001010100101001110001100110000;
		b = 32'b01010010000010111100101101110111;
		correct = 32'b00111000000010000101001101010100;
		#400 //4878744.0 * 150103500000.0 = 3.2502532e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011010000101100010101000001010;
		b = 32'b10111001111110101110001110111001;
		correct = 32'b00011111100110010011100100010100;
		#400 //-3.1053232e-23 * -0.00047853382 = 6.489245e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100110011011111011110011100010;
		b = 32'b10101101111100111000010110101000;
		correct = 32'b11110111111111000000010110010110;
		#400 //2.8303247e+23 * -2.7685257e-11 = -1.02232196e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010001011111011001110000101;
		b = 32'b11011001011110010000110010110100;
		correct = 32'b00100000001101001001101011001010;
		#400 //-0.0006702471 * -4381327300000000.0 = 1.5297808e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101010000100111011010110011111;
		b = 32'b01000101010001000110101110110111;
		correct = 32'b01100100010000001000001101101100;
		#400 //4.4642444e+25 * 3142.7322 = 1.4204979e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100110111110101111000001100010;
		b = 32'b01000111011011110101001100010000;
		correct = 32'b10011111000001100011011000111111;
		#400 //-1.7412391e-15 * 61267.062 = -2.8420475e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100001011101110001110100000001;
		b = 32'b11010111010111110011111011011010;
		correct = 32'b00001001100011011010111101010001;
		#400 //-8.372524e-19 * -245461040000000.0 = 3.4109382e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110111101100001011111101011011;
		b = 32'b11000111000000000101111010100100;
		correct = 32'b01110000001100000011110100001100;
		#400 //-7.1697297e+33 * -32862.64 = 2.1817265e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100100010011000110001011111100;
		b = 32'b00110001110010101001111010101111;
		correct = 32'b11110010000000010001110110111011;
		#400 //-1.5081073e+22 * 5.897014e-09 = -2.5574085e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110110010000011000000011100;
		b = 32'b01011000100011001000011001100000;
		correct = 32'b10011101101101100101100001100101;
		#400 //-5.966065e-06 * 1236070100000000.0 = -4.8266397e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110010100111100100100101111100;
		b = 32'b11011100101011010010100011000111;
		correct = 32'b11010101011010100000001101000101;
		#400 //6.270396e+30 * -3.8992005e+17 = -16081235000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100000101111111011100000110010;
		b = 32'b00110110001110111101111000000111;
		correct = 32'b10101010000000101001111111101000;
		#400 //-3.247855e-19 * 2.7994408e-06 = -1.1601798e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000011111101001101001100100001;
		b = 32'b10111001001010000001000100101001;
		correct = 32'b11001010001110100111010101101111;
		#400 //489.64944 * -0.00016028121 = -3054939.8
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100000111111110100001100000001;
		b = 32'b00110011100001100011111111001111;
		correct = 32'b11101100111100110110000100100000;
		#400 //-1.4714837e+20 * 6.251468e-08 = -2.353821e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011101110110100011011110100000;
		b = 32'b11011010101111001100111010010100;
		correct = 32'b00000010100100111111000001000000;
		#400 //-5.7761634e-21 * -2.6572215e+16 = 2.1737605e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110010010110001001101011011110;
		b = 32'b01110110111010001100010110010111;
		correct = 32'b00111010111011100011100001000111;
		#400 //4.290303e+30 * 2.3605869e+33 = 0.0018174731
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110110100100100100101111010010;
		b = 32'b00000101011110111110110011010110;
		correct = 32'b01110000100101001010100110011001;
		#400 //4.3599657e-06 * 1.1845463e-35 = 3.680705e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100110101111110100111011111111;
		b = 32'b01000001011011011001001100100110;
		correct = 32'b11100100110011100010010101000101;
		#400 //-4.517146e+23 * 14.848425 = -3.0421719e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010101010110100011010110101000;
		b = 32'b01111011100101111101010010110011;
		correct = 32'b00011001001101111111010111001101;
		#400 //14995249000000.0 * 1.5767018e+36 = 9.510517e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010011101111100100000011100011;
		b = 32'b01000011001110000111001011001100;
		correct = 32'b11010000000001000000011101001010;
		#400 //-1634264800000.0 * 184.44843 = -8860281000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010010101101100011110111001011;
		b = 32'b00110001000010001101100010100010;
		correct = 32'b01100001001010100111010111101101;
		#400 //391360380000.0 * 1.9913746e-09 = 1.9652775e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101011001001000011010010111011;
		b = 32'b10011001110100011000010001111101;
		correct = 32'b01010000110010001010001011001000;
		#400 //-5.833768e-13 * -2.1663605e-23 = 26928890000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111110111110100111101011000010;
		b = 32'b10110110001110100100010101110001;
		correct = 32'b01001000001011000001111100111011;
		#400 //-0.48921782 * -2.775658e-06 = 176252.92
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101100001011011100001101111001;
		b = 32'b10011110111000111111010110101100;
		correct = 32'b11001100110000110010001100110010;
		#400 //2.4693288e-12 * -2.4136167e-20 = -102308240.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100111011111000010100110001011;
		b = 32'b01111110011001011000000011111010;
		correct = 32'b00101000100011001010001100011111;
		#400 //1.1908027e+24 * 7.6265724e+37 = 1.5613865e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100111000011111001111111011000;
		b = 32'b00110001111010001111100100111100;
		correct = 32'b10110100100111011101000111011111;
		#400 //-1.9931888e-15 * 6.7804233e-09 = -2.939623e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001110000011000111101001101011;
		b = 32'b01010001000001001110100001110000;
		correct = 32'b00111100100001110100101001101010;
		#400 //589208260.0 * 35677210000.0 = 0.016514976
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110010101111110101000101110110;
		b = 32'b01100100100110001011110100001110;
		correct = 32'b10001101101000000101010011000011;
		#400 //-2.227237e-08 * 2.2540223e+22 = -9.881167e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110011100111111110011001101100;
		b = 32'b11011000010100011100011110100111;
		correct = 32'b10011010110000110010000101011110;
		#400 //7.445928e-08 * -922621700000000.0 = -8.070402e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001000110011100010000110001010;
		b = 32'b10010010001000000110100101110010;
		correct = 32'b00110110001001000111101100111100;
		#400 //-1.2406059e-33 * -5.061707e-28 = 2.4509636e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100101111000011100010111111010;
		b = 32'b11111011111000010110110101111100;
		correct = 32'b10101001100000000011001000111111;
		#400 //1.3327306e+23 * -2.3409748e+36 = -5.693058e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010110010011110000011101111111;
		b = 32'b10100010110101101010001111010111;
		correct = 32'b10110010111101101110110000111000;
		#400 //1.6723692e-25 * -5.817829e-18 = -2.8745589e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101010101111011101101100001101;
		b = 32'b10101101101000110110101110011000;
		correct = 32'b10111100100101001011010010101000;
		#400 //3.372514e-13 * -1.8578736e-11 = -0.01815255
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001011011010101111110001010001;
		b = 32'b00011110110101010111000011001000;
		correct = 32'b00101100000011001110101110101001;
		#400 //4.5256582e-32 * 2.2598897e-20 = 2.0026014e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001000011101110000100000010000;
		b = 32'b01001000101101001011000111010101;
		correct = 32'b00111111001011101111110111010100;
		#400 //252960.25 * 370062.66 = 0.6835606
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010111011000001011011101110100;
		b = 32'b11111110110110101001011011110000;
		correct = 32'b00011000000000111001011001111011;
		#400 //-247078530000000.0 * -1.4527771e+38 = 1.7007326e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110010010111011001011000000001;
		b = 32'b01100000000111101111001000011110;
		correct = 32'b00010001101100100111000111001100;
		#400 //1.2898e-08 * 4.5813e+19 = 2.815358e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101010001010101111011100111010;
		b = 32'b00110101101011010011110011100010;
		correct = 32'b11110011111111001010010001110111;
		#400 //-5.167122e+25 * 1.2907224e-06 = -4.0032793e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010110100110000111011100101;
		b = 32'b10101111001001111010010100111101;
		correct = 32'b01001011001000010010010101110100;
		#400 //-0.0016102461 * -1.5247266e-10 = 10560884.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001010100000110010001101111111;
		b = 32'b10101100011110011111111110111111;
		correct = 32'b01011101100001100100100101011001;
		#400 //-4297151.5 * -3.5526996e-12 = 1.2095454e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100100110010101100011011111100;
		b = 32'b10011000111100101001111110111010;
		correct = 32'b11001011010101011111010011100010;
		#400 //8.794063e-17 * -6.2716816e-24 = -14021858.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111101100100001001010100110;
		b = 32'b10111111000101000011101100111111;
		correct = 32'b11001000000110011100010010111100;
		#400 //91173.3 * -0.579029 = -157458.94
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001111100011101010010000110110;
		b = 32'b01010000100110101010110110100001;
		correct = 32'b10111110011011000001010000011011;
		#400 //-4786253000.0 * 20760562000.0 = -0.23054545
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111010010110001110001010111100;
		b = 32'b10111010001001010011100101110010;
		correct = 32'b10111111101010000000010110101111;
		#400 //0.0008273532 * -0.00063028105 = -1.3126734
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111111001110010010100110011000;
		b = 32'b00110011111110110011111010110111;
		correct = 32'b11001010101111001010101010110101;
		#400 //-0.7232909 * 1.1699506e-07 = -6182234.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011000101111011101101011010;
		b = 32'b10110110001101111000011110000101;
		correct = 32'b01010100010100111010010110000010;
		#400 //-9943898.0 * -2.7348008e-06 = 3636059400000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011110110110011101110101011111;
		b = 32'b11001000111101101101100101110100;
		correct = 32'b11010101011000011111000011011100;
		#400 //7.849404e+18 * -505547.62 = -15526537000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000100000010001110111011111010;
		b = 32'b00011011010001110000000011010101;
		correct = 32'b00101000001100000010011100011101;
		#400 //1.6096456e-36 * 1.6461163e-22 = 9.778444e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110110011110110010111011110001;
		b = 32'b10100000110111000011111011011001;
		correct = 32'b11010101000100011111101011101011;
		#400 //3.7429238e-06 * -3.731104e-19 = -10031679000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000100011101111001011011111110;
		b = 32'b11010011000110001011000110100111;
		correct = 32'b00110000110011111000110010010011;
		#400 //-990.35925 * -655815540000.0 = 1.5101186e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001011000100100001010111100100;
		b = 32'b11110101100100011001111000110100;
		correct = 32'b10010101000000000110100100110101;
		#400 //9573860.0 * -3.6918544e+32 = -2.5932388e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001111011101100110111010010000;
		b = 32'b00100101101110110010110011011110;
		correct = 32'b11101001001010001000010111010000;
		#400 //-4134441000.0 * 3.2469732e-16 = -1.2733216e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000011001011001111001111011111;
		b = 32'b00011101011100010011100000000011;
		correct = 32'b10100101001101111000110011111001;
		#400 //-5.0826207e-37 * 3.1925042e-21 = -1.5920483e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001100111100001010000011110010;
		b = 32'b10101000001100001010001100010011;
		correct = 32'b00100100001011100101111100011111;
		#400 //-3.707472e-31 * -9.805324e-15 = 3.7810806e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110101111001010111111011011111;
		b = 32'b00000101011001011110100000111001;
		correct = 32'b11101111111111111000101010110001;
		#400 //-1.7098754e-06 * 1.0810181e-35 = -1.5817269e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010010110010101010001000100000;
		b = 32'b00111010000011010010100111011100;
		correct = 32'b01011000001101111011110011011011;
		#400 //435151700000.0 * 0.00053849607 = 808087000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110001100001010000001011101111;
		b = 32'b10111110010101001001011010100000;
		correct = 32'b10110010101000000010110001001110;
		#400 //3.871143e-09 * -0.20760584 = -1.8646599e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100101011101011010001100000000;
		b = 32'b00011110000100010111000011111010;
		correct = 32'b01000110110110000010111000010011;
		#400 //2.1305589e-16 * 7.699599e-21 = 27671.037
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001010000010111111100101111010;
		b = 32'b10010110100001000100100101110011;
		correct = 32'b01110011000001110111000001000000;
		#400 //-2293342.5 * -2.1372103e-25 = 1.0730542e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101000011001010010100100001101;
		b = 32'b10110111111000100011110110110011;
		correct = 32'b00110000000000011010011011010100;
		#400 //-1.2720955e-14 * -2.697003e-05 = 4.7167004e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010100001111011000101001010010;
		b = 32'b10111001011010000010011101100010;
		correct = 32'b10011010010100010000001001100100;
		#400 //9.56934e-27 * -0.00022139915 = -4.3222118e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111111100110111111011011001111;
		b = 32'b01100000000001110110001100110010;
		correct = 32'b00011111000100110111010000101111;
		#400 //1.2184695 * 3.9022785e+19 = 3.1224566e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011110000010111111010000000111;
		b = 32'b10110011010111001001010010110010;
		correct = 32'b10101010001000100110110100000100;
		#400 //7.409062e-21 * -5.135798e-08 = -1.4426313e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011110010111001010101100000001;
		b = 32'b00111101001110101011110100111010;
		correct = 32'b01100000100101110100000110100110;
		#400 //3.975201e+18 * 0.045590617 = 8.71934e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100000111101101100001010011110;
		b = 32'b01100110111000110101000000010011;
		correct = 32'b10111001100010101111001101101100;
		#400 //-1.4224758e+20 * 5.3672715e+23 = -0.00026502775
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100111001101100101010100010011;
		b = 32'b01001111110101001110001100000110;
		correct = 32'b01010110110110110100000111111001;
		#400 //8.6104004e+23 * 7143296000.0 = 120538200000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000100011111100000111011100100;
		b = 32'b00111001000101100110000010001000;
		correct = 32'b00001010110110000100000010110000;
		#400 //2.9864394e-36 * 0.00014341075 = 2.0824376e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000101000000001011011110000011;
		b = 32'b00011001001101000101011001000111;
		correct = 32'b00101011001101101011100011001010;
		#400 //6.052237e-36 * 9.3232055e-24 = 6.4915835e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001110110000001000001011010101;
		b = 32'b10101100111101110101000111101010;
		correct = 32'b01100001010001110100010001111010;
		#400 //-1614899800.0 * -7.0292565e-12 = 2.2973977e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010001000010000101111010111000;
		b = 32'b11100111110001010001110100010100;
		correct = 32'b00101000101100010001110000010010;
		#400 //-36606540000.0 * -1.8616852e+24 = 1.9663121e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100001101011000000000001110000;
		b = 32'b00111011001001101011010111100100;
		correct = 32'b10100110000001000001000000000101;
		#400 //-1.1655289e-18 * 0.0025438005 = -4.581841e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100110101111110101101101001110;
		b = 32'b01111101011011101101110100101011;
		correct = 32'b10101000110011010001010110100110;
		#400 //-4.5182814e+23 * 1.984404e+37 = -2.276896e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011010111100000010001100000101;
		b = 32'b10100000010001000111001001010110;
		correct = 32'b11111010000111000111011110101101;
		#400 //3.379625e+16 * -1.6639676e-19 = -2.031064e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000101101101011010110001000001;
		b = 32'b00011101100101010101110010000001;
		correct = 32'b00100111100110111011000010111110;
		#400 //1.7084434e-35 * 3.953562e-21 = 4.3212766e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111001100010111100111011111111;
		b = 32'b11010000111110011011000101000111;
		correct = 32'b01101000000011110101011100011110;
		#400 //-9.074096e+34 * -33513159000.0 = 2.7076217e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001000101101000010010011101110;
		b = 32'b00000001111111000100000110111011;
		correct = 32'b11000110001101101101000101000010;
		#400 //-1.0842038e-33 * 9.26645e-38 = -11700.314
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111101011110101000001011111010;
		b = 32'b10110100001101111100111101100100;
		correct = 32'b11001000101011100111001011110000;
		#400 //0.061160065 * -1.7118651e-07 = -357271.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100101100000110001100111001001;
		b = 32'b01110010111000110001001000111010;
		correct = 32'b00110010000100111100110110001100;
		#400 //7.738821e+22 * 8.995217e+30 = 8.603262e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000111100011001011010100101110;
		b = 32'b10100101001001000001001000101101;
		correct = 32'b00100001110110111000101111011010;
		#400 //-2.1171347e-34 * -1.4230891e-16 = 1.4877036e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101011111110110111011001010011;
		b = 32'b11011111100011110111110111110000;
		correct = 32'b11001011111000000101000000111001;
		#400 //6.079983e+26 * -2.0679368e+19 = -29401202.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110110111000101000001100100100;
		b = 32'b01111100011101011110010010100011;
		correct = 32'b10111001111010111101001010010011;
		#400 //-2.2971073e+33 * 5.107e+36 = -0.00044979583
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011001010110000001001101000100;
		b = 32'b01101011100100111011101001000110;
		correct = 32'b10101101001110110011100001101111;
		#400 //-3801236000000000.0 * 3.571835e+26 = -1.064225e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001100111000100101100000110100;
		b = 32'b10011110101001110010001001110010;
		correct = 32'b11101101101011010101100010010010;
		#400 //118669730.0 * -1.7696059e-20 = -6.7059977e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010000100101110101000010010010;
		b = 32'b00000000111110110101010011010100;
		correct = 32'b11001111000110100010000000100000;
		#400 //-5.9683137e-29 * 2.308114e-38 = -2585796600.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101010111111101001110111101111;
		b = 32'b01000111000100100110101001111011;
		correct = 32'b01100011010111101001011101110111;
		#400 //1.5390649e+26 * 37482.48 = 4.1060914e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001000001011000101010101100011;
		b = 32'b00001011010011100101000101101111;
		correct = 32'b11111100010101011101010011110110;
		#400 //-176469.55 * 3.973542e-32 = -4.4411144e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000010111100000110000000011011;
		b = 32'b00100111110000110000100101110110;
		correct = 32'b00011010100111011100000101000111;
		#400 //3.5319992e-37 * 5.413363e-15 = 6.5245934e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101000000011010011110001001111;
		b = 32'b11110001010000000010000111011101;
		correct = 32'b10110110001111000010111100111001;
		#400 //2.6678647e+24 * -9.5139296e+29 = -2.804167e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000111111010010100101001001100;
		b = 32'b01110001100111111010000111000100;
		correct = 32'b10010101101110110001000000000011;
		#400 //-119444.59 * 1.5809177e+30 = -7.555396e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010111101000010010010011010111;
		b = 32'b01001111000001100000110100001100;
		correct = 32'b11001000000110011101111010110111;
		#400 //-354359200000000.0 * 2249002000.0 = -157562.86
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010001101110100101010011011110;
		b = 32'b11010111001110000110001011110001;
		correct = 32'b10111010000000010101100110101000;
		#400 //100035970000.0 * -202735090000000.0 = -0.00049343193
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011111001110010100000010100100;
		b = 32'b11010110111110010001100010000011;
		correct = 32'b11000111101111100110001100011111;
		#400 //1.334885e+19 * -136941840000000.0 = -97478.24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011100111110000100010011001110;
		b = 32'b01010001000100000001000101101100;
		correct = 32'b10001011010111001001010001000000;
		#400 //-1.6429049e-21 * 38672974000.0 = -4.248199e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010111111100000101011110111;
		b = 32'b10110000001110110111111100101010;
		correct = 32'b01001010001011010110110111111010;
		#400 //-0.001938193 * -6.8210915e-10 = 2841470.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111111011100101100000100000111;
		b = 32'b10111001100100000101111110010001;
		correct = 32'b11000101010101110011100100110001;
		#400 //0.94825786 * -0.00027537023 = -3443.5745
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101001001011000101001100111100;
		b = 32'b00101011111100111100111011111110;
		correct = 32'b00111100101101001111000100101110;
		#400 //3.8263866e-14 * 1.732364e-12 = 0.02208766
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100111100010100111110100111101;
		b = 32'b10011000010101000011101010101001;
		correct = 32'b01001110101001110000110100111100;
		#400 //-3.843848e-15 * -2.7429974e-24 = 1401331200.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101011100011110111001001110101;
		b = 32'b10010001101110111110110001110101;
		correct = 32'b01011001010000110110100101011100;
		#400 //-1.0192529e-12 * -2.9649126e-28 = 3437716500000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000011110111010001111101110100;
		b = 32'b01011011110011000110001000001010;
		correct = 32'b00100111100010100111101111011001;
		#400 //442.24573 * 1.1505738e+17 = 3.843697e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110110100101001110100000000100;
		b = 32'b10111101100101110010101010001100;
		correct = 32'b01111000011111000010110001000010;
		#400 //-1.5100894e+33 * -0.07381162 = 2.0458695e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111011010010001111001111111011;
		b = 32'b01000000010110100011100000101111;
		correct = 32'b10111010011010111011111010000110;
		#400 //-0.0030663002 * 3.4096792 = -0.0008992929
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100011101001010110100111110111;
		b = 32'b10101100100111110000001011011001;
		correct = 32'b11110110100001010010011101110011;
		#400 //6.1026967e+21 * -4.519368e-12 = -1.350343e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101101111110011111110010010001;
		b = 32'b00101110100101001001100000010110;
		correct = 32'b11111110110101110101011100011001;
		#400 //-9.6708877e+27 * 6.757277e-11 = -1.4311813e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100000101100011001110000001011;
		b = 32'b10100010110100110100110011000010;
		correct = 32'b00111101010101110010111010111101;
		#400 //-3.0088227e-19 * -5.7272935e-18 = 0.052534807
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000000101010110010100001011100;
		b = 32'b00000100010101110000110101111101;
		correct = 32'b11111011110010111011111101000001;
		#400 //-5.3486767 * 2.5279322e-36 = -2.1158307e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100001010101001010001010111011;
		b = 32'b11011111110111110101000011111110;
		correct = 32'b01000000111100111100000110010000;
		#400 //-2.4515223e+20 * -3.2183281e+19 = 7.617378
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110000010000101011010011011000;
		b = 32'b10010001110110011110010001101000;
		correct = 32'b11011101111001001100001001011010;
		#400 //7.0833783e-10 * -3.437733e-28 = -2.0604796e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011110011001111000111100001110;
		b = 32'b10101110011100000100100100101111;
		correct = 32'b11101111011101101011001111000100;
		#400 //4.1713926e+18 * -5.4634682e-11 = -7.6350636e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111111010010101110010110111101;
		b = 32'b11110110101110000100111011010001;
		correct = 32'b10001000000011001110100100000110;
		#400 //0.792568 * -1.869104e+33 = -4.2403635e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111010011100100101010011111011;
		b = 32'b10011100000000000000100010110000;
		correct = 32'b11011101111100100100010010001010;
		#400 //0.00092442305 * -4.2362876e-22 = -2.1821537e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100111111100000010110110100101;
		b = 32'b11010101011110111001011101001101;
		correct = 32'b10010001111101000110001100100101;
		#400 //6.666287e-15 * -17289203000000.0 = -3.8557515e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000100000111100001000010010110;
		b = 32'b11000000101000100101010000001000;
		correct = 32'b10000010111110010100011010111100;
		#400 //1.8580427e-36 * -5.0727577 = -3.6627861e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111000001111101100100001010001;
		b = 32'b11011011100001111001010110100100;
		correct = 32'b11011100001101000001110000110110;
		#400 //1.5478114e+34 * -7.632731e+16 = -2.0278606e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010000001100101011000101111010;
		b = 32'b10000010110011010010111101010110;
		correct = 32'b01001100110111101111001010010100;
		#400 //-3.5241033e-29 * -3.0149212e-37 = 116888740.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111110000110011011110000001101;
		b = 32'b10000001010001000111001000000101;
		correct = 32'b01111100010010000101011101000111;
		#400 //-0.15013142 * -3.608132e-38 = 4.1609183e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100100010011001010110110100011;
		b = 32'b01010111110001111101100000011010;
		correct = 32'b00001100000000110001100010100100;
		#400 //4.4382525e-17 * 439461930000000.0 = 1.0099288e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001101111000000101111110010000;
		b = 32'b11001110001111000111010111110010;
		correct = 32'b00111111000110000110010000101111;
		#400 //-470544900.0 * -790461600.0 = 0.5952787
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010110100101001110010001011110;
		b = 32'b00111100111001111001000101101110;
		correct = 32'b00011001001001001001100111100011;
		#400 //2.405481e-25 * 0.028267588 = 8.5096785e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110001110111010010100001111001;
		b = 32'b00111000101101100010011011000001;
		correct = 32'b10111000100110110110100100010110;
		#400 //-6.4365477e-09 * 8.685655e-05 = -7.41055e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111100111100011010100101101110;
		b = 32'b00011011011101001111110101010001;
		correct = 32'b11100000111111001000010111010100;
		#400 //-0.029499736 * 2.0265058e-22 = -1.4556946e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110101000011011001100011000001;
		b = 32'b01101101000000111011101010111111;
		correct = 32'b00000111100010011001011001111110;
		#400 //5.274888e-07 * 2.5480187e+27 = 2.070192e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101100100001011000111101010101;
		b = 32'b10011101000111111010100010010001;
		correct = 32'b11001110110101100010011100101000;
		#400 //3.7960004e-12 * -2.1130622e-21 = -1796445200.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101001110110011101001001001001;
		b = 32'b11001110110011000110010101101011;
		correct = 32'b11011010100010000110100001001001;
		#400 //3.2916243e+25 * -1714599300.0 = -1.919763e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001000000001010101000000010101;
		b = 32'b01000100000010010100000100100000;
		correct = 32'b01000011011110001010010111111100;
		#400 //136512.33 * 549.0176 = 248.64838
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101101110111100000111111001100;
		b = 32'b10111000110000000110001011001011;
		correct = 32'b01110100100100111011111010000011;
		#400 //-8.590596e+27 * -9.173675e-05 = 9.3644e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111101000111110111110001100110;
		b = 32'b00000010101110100011001011100111;
		correct = 32'b11111001110110110100010111101011;
		#400 //-0.038936995 * 2.735946e-37 = -1.4231639e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111000001010001011101001100100;
		b = 32'b00000011111011100000110000001110;
		correct = 32'b01110011101101010111010000000001;
		#400 //4.022791e-05 * 1.399115e-36 = 2.8752398e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110110010000101100100101011010;
		b = 32'b01001011111010010100100110111001;
		correct = 32'b01101001110101011100000000001101;
		#400 //9.8768504e+32 * 30577522.0 = 3.2301017e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111011100001001100011011111100;
		b = 32'b11101000100101011101010001010010;
		correct = 32'b10010010011000101101110101011000;
		#400 //0.004052041 * -5.660394e+24 = -7.1585853e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011001011000011100010010111101;
		b = 32'b10111011010111101011011011101110;
		correct = 32'b01011101100000011100000101010100;
		#400 //-3971761600000000.0 * -0.0033983546 = 1.1687308e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111010111011001100100100111001;
		b = 32'b01010010001100011000000000111000;
		correct = 32'b00101000001010101100000001111110;
		#400 //0.001806534 * 190590090000.0 = 9.478636e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101010011101101110110001000000;
		b = 32'b10000000000011110001010011000011;
		correct = 32'b11101011000000101111101111100111;
		#400 //2.1931155e-13 * -1.38498e-39 = -1.5834993e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100100110011001000000101110011;
		b = 32'b00101001110010010110010010011101;
		correct = 32'b00111010100000011111101001110011;
		#400 //8.869019e-17 * 8.943647e-14 = 0.0009916559
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111000101011101000011011100000;
		b = 32'b10010010111100110000100011101011;
		correct = 32'b01100101001101111101011001011011;
		#400 //-8.322089e-05 * -1.5337654e-27 = 5.42592e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010001111001000000010010100111;
		b = 32'b10010001001111101100011111011010;
		correct = 32'b01000000000110001111101111010001;
		#400 //-3.5974925e-28 * -1.5049941e-28 = 2.3903697
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110010011110110110100101011110;
		b = 32'b10001111011101110100111111001001;
		correct = 32'b11100010100000100001111100111010;
		#400 //1.4634081e-08 * -1.2193406e-29 = -1.2001634e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011110100010001011110010001110;
		b = 32'b00111111111110111100110011001000;
		correct = 32'b00011110000010110000010001110000;
		#400 //1.4477544e-20 * 1.9671869 = 7.359516e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010001000010100110001000001011;
		b = 32'b11111010110101100011011011010101;
		correct = 32'b00010101101001010110000001110010;
		#400 //-37146900000.0 * -5.5613183e+35 = 6.6795133e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110101001111001110111000101011;
		b = 32'b00101100110011010010011000110001;
		correct = 32'b11000111111010111100001011001110;
		#400 //-7.038204e-07 * 5.8306905e-12 = -120709.61
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111010011010010011010101010110;
		b = 32'b01111110010000010000101100011001;
		correct = 32'b00111011100110101010000111000111;
		#400 //3.0272174e+35 * 6.4149656e+37 = 0.0047189924
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101000110101001001100011110001;
		b = 32'b00101000101110101001111100000011;
		correct = 32'b00111111100100011101000100010000;
		#400 //2.3603056e-14 * 2.0719109e-14 = 1.1391926
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111000100011011110111000011000;
		b = 32'b01010011111011010011101111001111;
		correct = 32'b00100100000110010010100001001110;
		#400 //6.767752e-05 * 2037821300000.0 = 3.3210726e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101011001010101100100011011101;
		b = 32'b01011000101001001011110110010011;
		correct = 32'b10010010000001001011001000110110;
		#400 //-6.0674886e-13 * 1449073000000000.0 = -4.187152e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110000111011000110011110001;
		b = 32'b00010100100001011101101000110111;
		correct = 32'b11100001000101101010100101111001;
		#400 //-2.3476862e-06 * 1.3515639e-26 = -1.7370146e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100110111100001010110001110000;
		b = 32'b10110101011100111111111101101111;
		correct = 32'b01110000111111001000001100100101;
		#400 //-5.6827443e+23 * -9.089626e-07 = 6.2519013e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110000011011001001001001110010;
		b = 32'b01100010100000111110110100111111;
		correct = 32'b01001101011001011000011111010101;
		#400 //2.9286202e+29 * 1.2168094e+21 = 240680270.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000111110110111010010110000001;
		b = 32'b00000111010001100111000100010101;
		correct = 32'b11000000000011011010110101111001;
		#400 //-3.3048732e-34 * 1.4929096e-34 = -2.213713
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010111011001110010001101010000;
		b = 32'b10001011001010111001010101101100;
		correct = 32'b01001011101011000110110101001111;
		#400 //-7.4684696e-25 * -3.3045815e-32 = 22600350.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101011101100101111111011001110;
		b = 32'b01011110011111001110010110001000;
		correct = 32'b11001100101101010011000100011101;
		#400 //-4.3278415e+26 * 4.5557803e+18 = -94996710.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111110001000111000111000001001;
		b = 32'b11000101101110110101101010001111;
		correct = 32'b00110111110111110111101100101110;
		#400 //-0.15972151 * -5995.32 = 2.6641032e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011001110110100011011110100001;
		b = 32'b00001001100110110011110111010111;
		correct = 32'b11001111101100111110110011000011;
		#400 //-2.256314e-23 * 3.7373047e-33 = -6037276000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110011110000011000010010111000;
		b = 32'b01101010001100100100100010110001;
		correct = 32'b01001001000010101111000000001100;
		#400 //3.066422e+31 * 5.388302e+25 = 569088.75
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111011101000000000001101011001;
		b = 32'b00111100110100001001011001100110;
		correct = 32'b00111110010001000110001001101110;
		#400 //0.0048832116 * 0.02546234 = 0.19178173
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110110000010011111001100010100;
		b = 32'b11110100000001101101111000001110;
		correct = 32'b10000001100000101110110011011001;
		#400 //2.055608e-06 * -4.2741185e+31 = -4.809432e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001010000001110010101110101000;
		b = 32'b01100010010010110011001101001001;
		correct = 32'b10100111001010100100101100010110;
		#400 //-2214634.0 * 9.370961e+20 = -2.3632943e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001101010011100000101010111111;
		b = 32'b01001000010010101000110101000011;
		correct = 32'b00000100100000100011010010100000;
		#400 //6.3491586e-31 * 207413.05 = 3.061118e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010000000101111010000011100111;
		b = 32'b11100110110010010001001000101010;
		correct = 32'b10101000110000010000110011111111;
		#400 //10175618000.0 * -4.7476537e+23 = -2.143294e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100111011001110000010100010111;
		b = 32'b01101100010011010010111101000010;
		correct = 32'b00111010100100000001110111100110;
		#400 //1.09096055e+24 * 9.9221185e+26 = 0.0010995239
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100110010100001101010111010000;
		b = 32'b00110100011101110101000101010101;
		correct = 32'b10110001010110000010101010100010;
		#400 //-7.2454267e-16 * 2.3033256e-07 = -3.145637e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111110000010010011010100001011;
		b = 32'b11111100111001110011101100000100;
		correct = 32'b01000000100101111110011110100101;
		#400 //-4.5594913e+37 * -9.6049404e+36 = 4.747027
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011001110100011001110101010001;
		b = 32'b01110011011101110111110110010001;
		correct = 32'b00100101110110001101001001011101;
		#400 //7375155000000000.0 * 1.9608217e+31 = 3.7612575e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001001000000001010000000100010;
		b = 32'b11000111000011111111010010011010;
		correct = 32'b00000001011001001011110100000010;
		#400 //-1.5482734e-33 * -36852.6 = 4.2012593e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111000101011100101100101101;
		b = 32'b01001100011010110111001001010100;
		correct = 32'b00111010001000101101111010110101;
		#400 //38347.176 * 61720910.0 = 0.00062129955
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010101001101101001001100100110;
		b = 32'b01001100101111011101100111011000;
		correct = 32'b00000111111101100011000001001011;
		#400 //3.6870687e-26 * 99536580.0 = 3.704235e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111110100111110000101100101;
		b = 32'b01010101000001100011110110000111;
		correct = 32'b00110010010010100000011111101001;
		#400 //108482.79 * 9224926000000.0 = 1.1759746e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111011100010011000001010111100;
		b = 32'b00001001010100010000011110000100;
		correct = 32'b11110001101010000110100100010101;
		#400 //-0.004196493 * 2.5160994e-33 = -1.6678566e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111000000100001000101111010;
		b = 32'b11100111100001000110001111011001;
		correct = 32'b00001110111110111000001010101101;
		#400 //-7.752673e-06 * -1.2503885e+24 = 6.2002113e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001101010001110010100000011001;
		b = 32'b00000111110011100111101000011110;
		correct = 32'b11000100111101101110110010000000;
		#400 //-6.1369875e-31 * 3.106721e-34 = -1975.3906
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010111101000010101011111110001;
		b = 32'b11001111110101001010111010010000;
		correct = 32'b10000111010000100011010010001100;
		#400 //1.0426581e-24 * -7136420000.0 = -1.461038e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011110101011100011110000011100;
		b = 32'b00100100001000100010100101010110;
		correct = 32'b11111010000010011000011110101001;
		#400 //-6.2774703e+18 * 3.5163163e-17 = -1.7852405e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001010110000100101111001110000;
		b = 32'b00011011110101101011011111011001;
		correct = 32'b11101110011001111011110100000111;
		#400 //-6369080.0 * 3.552214e-22 = -1.7929889e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001000110000101001001100100111;
		b = 32'b00101100011001100001111011000001;
		correct = 32'b10011011110110000111010100001001;
		#400 //-1.1710546e-33 * 3.2702038e-12 = -3.5809835e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011001001110000111110111000100;
		b = 32'b10010101111101001010011010111111;
		correct = 32'b11000010110000010000110010011101;
		#400 //9.537975e-24 * -9.8813894e-26 = -96.524635
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011011101100101000100101000001;
		b = 32'b01000010110000100011101001101100;
		correct = 32'b01011000011010110101000100111001;
		#400 //1.0050692e+17 * 97.114105 = 1034936300000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001111111110111001010101011001;
		b = 32'b00111101110000111100101011110011;
		correct = 32'b01010001101001000111100100100111;
		#400 //8441737700.0 * 0.09560194 = 88300904000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000000000111001001010011110100;
		b = 32'b10111010110000111100000010011010;
		correct = 32'b00000100000101011000001110110110;
		#400 //-2.624828e-39 * -0.0014934719 = 1.7575345e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101001100100011110111110011000;
		b = 32'b11100110011001000011100000100101;
		correct = 32'b10000010101000111011001101001110;
		#400 //6.4808564e-14 * -2.6943381e+23 = -2.4053613e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100010110011110001001011101110;
		b = 32'b01100010010010000100010000110111;
		correct = 32'b01000000000001000101100111011010;
		#400 //1.90992e+21 * 9.2356605e+20 = 2.067984
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111110110000011100110010000100;
		b = 32'b01011110111110100110010110101101;
		correct = 32'b01011111010001100010001010100010;
		#400 //1.2880145e+38 * 9.021509e+18 = 1.4277152e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000100010101011101110101011100;
		b = 32'b00000001011110101111000111111001;
		correct = 32'b01000010010110100010110000101101;
		#400 //2.5139673e-36 * 4.6091355e-38 = 54.54314
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000000110111011001001011100011;
		b = 32'b10101001010100100101010010001000;
		correct = 32'b01010111000001101101011110101100;
		#400 //-6.9241805 * -4.6702686e-14 = 148260860000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111110011111101111110101010110;
		b = 32'b01100001011010000011000100111011;
		correct = 32'b11011100100011001001000101000001;
		#400 //-8.4734827e+37 * 2.676995e+20 = -3.1652964e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100110010101101011101001111100;
		b = 32'b00010011111000100110001001111111;
		correct = 32'b11010001111100101101000110100000;
		#400 //-7.44989e-16 * 5.7147545e-27 = -130362380000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111011010100111100001001011010;
		b = 32'b01101111010000001111010110010111;
		correct = 32'b11001011100011000111100010001110;
		#400 //-1.09951656e+36 * 5.971802e+28 = -18411804.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011001111111001101100111000110;
		b = 32'b01000100101011010011110001110101;
		correct = 32'b00010100101110101101001101000011;
		#400 //2.6144147e-23 * 1385.8893 = 1.8864528e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010010110110001010110111100100;
		b = 32'b11111000101011110011100011001111;
		correct = 32'b00011001100111100100100011100001;
		#400 //-465315170000.0 * -2.843138e+34 = 1.6366253e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101001011101001100001001000001;
		b = 32'b10011100101111111000101000100001;
		correct = 32'b01001100001000111001000010010101;
		#400 //-5.4347372e-14 * -1.2675025e-21 = 42877524.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001101111001010100100011100011;
		b = 32'b11010010110111110000101010110010;
		correct = 32'b00111010100000111001010100101101;
		#400 //-480844900.0 * -478978570000.0 = 0.0010038965
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100100001011101111000110110111;
		b = 32'b11000010100110100101010010001001;
		correct = 32'b10100001000100010001100011011000;
		#400 //3.7934976e-17 * -77.16511 = -4.916079e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010110110001111000110101000010;
		b = 32'b10100110100000111011101001111000;
		correct = 32'b11101111110000011110011101011100;
		#400 //109704760000000.0 * -9.140493e-16 = -1.2002061e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100101001010011010010011111110;
		b = 32'b01010110000110101110000101100100;
		correct = 32'b01001110100011000011001110100001;
		#400 //5.007022e+22 * 42573210000000.0 = 1176096900.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100111010111011000100011110011;
		b = 32'b11000111011001011101100101000001;
		correct = 32'b10011111011101101011110110001011;
		#400 //3.0744151e-15 * -58841.254 = -5.2249313e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111010111101101101010001111000;
		b = 32'b00011101101000010000000111010101;
		correct = 32'b01011100110001000011101010010000;
		#400 //0.0018831631 * 4.261824e-21 = 4.418679e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100010011010011110010011000001;
		b = 32'b11001011011010010101011000101010;
		correct = 32'b11010110100000000100111000111000;
		#400 //1.0786437e+21 * -15291946.0 = -70536720000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001100011001010111011001101111;
		b = 32'b00111110010000000011000010101001;
		correct = 32'b10001101100110001101001011100100;
		#400 //-1.7677158e-31 * 0.18768562 = -9.418493e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001111100100000001101110111001;
		b = 32'b10100100110000011011100101011111;
		correct = 32'b11101010001111100110111100110001;
		#400 //4835472000.0 * -8.401444e-17 = -5.755525e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111000011011000101100000010000;
		b = 32'b11010010100010001110111110000110;
		correct = 32'b11100101010111001110101111101010;
		#400 //1.9174503e+34 * -294067040000.0 = -6.520453e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111001100110000101011001000110;
		b = 32'b11011010001011000101001111011110;
		correct = 32'b00011110111000100100110110011001;
		#400 //-0.00029055978 * -1.2126477e+16 = 2.3960774e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111000101010110000011011001101;
		b = 32'b11001000101111000011000010101101;
		correct = 32'b11101111011010001010011011100101;
		#400 //2.7750647e+34 * -385413.4 = -7.2002285e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011100000110100110101111101010;
		b = 32'b10011100000110110111010001110011;
		correct = 32'b10111111011111100100110001011110;
		#400 //5.10938e-22 * -5.1435705e-22 = -0.9933528
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101110011000011100100111010101;
		b = 32'b11100100000000110000111101011100;
		correct = 32'b11001001110111001000010001000101;
		#400 //1.7469532e+28 * -9.670521e+21 = -1806472.6
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110111001101001011110010011010;
		b = 32'b10110111100000011001010010111011;
		correct = 32'b11111111001100101000100000011000;
		#400 //3.6657763e+33 * -1.5447256e-05 = -2.3730922e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000001100001010000100011100100;
		b = 32'b10000101001001001000111101001100;
		correct = 32'b11111011110011101111010100100101;
		#400 //16.629341 * -7.7375624e-36 = -2.1491705e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000000000110000000110010110111;
		b = 32'b00000111111110011101001000101010;
		correct = 32'b11110111100110111100111101111010;
		#400 //-2.375776 * 3.758888e-34 = -6.320423e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010101110111111001010101111101;
		b = 32'b11000011010001110001011110001110;
		correct = 32'b10010010000011111011111100001111;
		#400 //9.0304834e-26 * -199.09201 = -4.535834e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011101100111101010111011010101;
		b = 32'b00000100100001111100111100110100;
		correct = 32'b01011000100101011000111011101010;
		#400 //4.2003024e-21 * 3.1928633e-36 = 1315528400000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111101111011000101111000010001;
		b = 32'b11011000111100110100101001000100;
		correct = 32'b00100100011110001011011100111000;
		#400 //-0.11541379 * -2140002400000000.0 = 5.393162e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010100100000110011000000000010;
		b = 32'b00110000100100001000101010111101;
		correct = 32'b10100011011010000101100100001011;
		#400 //-1.3246555e-26 * 1.0516811e-09 = -1.2595601e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100011000011000110100011010010;
		b = 32'b10100000001001110100011100101111;
		correct = 32'b11000010010101101110000101110011;
		#400 //7.611612e-18 * -1.4169003e-19 = -53.720165
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100011100100111011111000110000;
		b = 32'b01111101001001011011011011000000;
		correct = 32'b10100101111001000011110011101000;
		#400 //-5.4507517e+21 * 1.376697e+37 = -3.9592967e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000000110001111001001111110000;
		b = 32'b10111011100111011100000000101110;
		correct = 32'b10000100101000011111000001011001;
		#400 //1.8328334e-38 * -0.0048141694 = -3.8071643e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000101100010000111101110011000;
		b = 32'b01000110000000111001001111110110;
		correct = 32'b00111111000001001100010101111101;
		#400 //4367.449 * 8420.99 = 0.51863843
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001100001011111101011110111011;
		b = 32'b00000111101001110101100001110011;
		correct = 32'b11000100000001100111111111010111;
		#400 //-1.3546429e-31 * 2.5179353e-34 = -537.9975
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001010000000110101111100011011;
		b = 32'b00100011111010000000100111110001;
		correct = 32'b11100101100100001110111111111010;
		#400 //-2152390.8 * 2.51577e-17 = -8.5555945e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001100101001100000101000110000;
		b = 32'b00011011111011101100110000011101;
		correct = 32'b11110000001100100000000001001001;
		#400 //-87052670.0 * 3.9505702e-22 = -2.203547e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001001010011001010101100111110;
		b = 32'b10110011111111100100101111111111;
		correct = 32'b11010100110011100000101000101000;
		#400 //838323.9 * -1.184162e-07 = -7079469000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100101100000101011111110000111;
		b = 32'b10010000001111100101111101001010;
		correct = 32'b01010100101011111101001001001101;
		#400 //-2.268119e-16 * -3.75443e-29 = 6041180300000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100111000001100101111011110000;
		b = 32'b10101110100010001101100110100111;
		correct = 32'b10110111111110110101110010101010;
		#400 //1.8647701e-15 * -6.223227e-11 = -2.9964682e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011010101011100010001111000001;
		b = 32'b01000010000111001101001101000001;
		correct = 32'b00011000000011100010000111001001;
		#400 //7.2022477e-23 * 39.206303 = 1.8370127e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010110000101110111010101000111;
		b = 32'b10111111010100101000011101000110;
		correct = 32'b00010110001110000010101111010110;
		#400 //-1.2234689e-25 * -0.8223766 = 1.4877234e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100101011001111011011111001000;
		b = 32'b11001001110011001100110010101001;
		correct = 32'b00011011000100001101001011110110;
		#400 //-2.0098324e-16 * -1677717.1 = 1.1979566e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001101111101001011011010100111;
		b = 32'b00000011000111000001011001001011;
		correct = 32'b01001010010010001010110110110100;
		#400 //1.5081633e-30 * 4.586987e-37 = 3287917.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110110011100101000100000001001;
		b = 32'b01010010010101101101001101011010;
		correct = 32'b11100011100100001000001000001101;
		#400 //-1.2297802e+33 * 230667220000.0 = -5.3314046e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010010011010000001100111111000;
		b = 32'b01111010000111111001001111111111;
		correct = 32'b00010111101110100010110000001100;
		#400 //249217020000.0 * 2.0714423e+35 = 1.2031087e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010101100111000111110000010000;
		b = 32'b11010110111000110010111011101100;
		correct = 32'b10111110001100000101010101101011;
		#400 //21507082000000.0 * -124895330000000.0 = -0.17220084
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001000110100001010011111001011;
		b = 32'b01100100111100111101010011101001;
		correct = 32'b10100011010110110001000101111100;
		#400 //-427326.34 * 3.5983205e+22 = -1.1875716e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110111101001110000011001000110;
		b = 32'b11011110001111100110010100110110;
		correct = 32'b01011000111000001001001110000101;
		#400 //-6.775319e+33 * -3.4298578e+18 = 1975393600000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011101000111111111010101011100;
		b = 32'b01001001100001011011111000001001;
		correct = 32'b11010011000110010001011100101011;
		#400 //-7.2038875e+17 * 1095617.1 = -657518700000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110100001011100101001000001110;
		b = 32'b01100100110100111100110101001100;
		correct = 32'b10001110110100101011001001110101;
		#400 //-1.6234864e-07 * 3.125645e+22 = -5.1940845e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110111100011010101011111100101;
		b = 32'b00110100001000011110100011101100;
		correct = 32'b01000010110111110111101101010011;
		#400 //1.6849439e-05 * 1.507903e-07 = 111.74087
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100001111110110101011100011000;
		b = 32'b10100110100111001101010100001001;
		correct = 32'b00111010110011010010001000110011;
		#400 //-1.7031475e-18 * -1.0882418e-15 = 0.0015650451
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110101110101111011011011101100;
		b = 32'b11101100101110000011000111101000;
		correct = 32'b10001000100101011110011101001010;
		#400 //1.6071986e-06 * -1.7814242e+27 = -9.021987e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101001000111100001010011100011;
		b = 32'b01111000110011001101111101100010;
		correct = 32'b00101111110001011000100000101111;
		#400 //1.1944307e+25 * 3.3242478e+34 = 3.5930856e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100011111010110001000010001011;
		b = 32'b11110110101010101101010111001110;
		correct = 32'b10101100101100000001111111100100;
		#400 //8.672354e+21 * -1.7324745e+33 = -5.0057614e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110100100000101101110001100011;
		b = 32'b01110000000001001001010110101010;
		correct = 32'b11000011111111001010101111110111;
		#400 //-8.294294e+31 * 1.6413182e+29 = -505.34348
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010110011100100010001101011111;
		b = 32'b11010010000100110110100000100011;
		correct = 32'b10000011110100100100001001110011;
		#400 //1.9559765e-25 * -158276830000.0 = -1.2357947e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101100101101110100110011001010;
		b = 32'b00010101000001000101100110000110;
		correct = 32'b01010111001100010100011010011001;
		#400 //5.209698e-12 * 2.672781e-26 = 194916770000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011111011110101100000011000100;
		b = 32'b00110000010011010111101101111100;
		correct = 32'b00101110100111000011001100111111;
		#400 //5.309901e-20 * 7.475405e-10 = 7.103162e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010110001000100011011000100101;
		b = 32'b10101001010011100100011101110101;
		correct = 32'b11101100010010010100111101111010;
		#400 //44588360000000.0 * -4.5803168e-14 = -9.734776e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000110011000110000111010010101;
		b = 32'b10000011011100110010101111101100;
		correct = 32'b11000010011011110000100100001000;
		#400 //4.2704668e-35 * -7.14617e-37 = -59.75882
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101011001110000001010011110000;
		b = 32'b01011100010111001100001111000100;
		correct = 32'b01001110010101010111011001011000;
		#400 //2.2254123e+26 * 2.4855897e+17 = 895325700.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100111011100010000110100100110;
		b = 32'b00111000001100011111110101111100;
		correct = 32'b11101110101011010101100110010001;
		#400 //-1.1383329e+24 * 4.2436164e-05 = -2.6824593e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110111001001101100000011100100;
		b = 32'b11010000000110001111011100101111;
		correct = 32'b11100110100010111000100110011111;
		#400 //3.3821624e+33 * -10265345000.0 = -3.294738e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010101010111000100101000111010;
		b = 32'b10011000001001011101110100000000;
		correct = 32'b11111100101010100000000010001100;
		#400 //15138210000000.0 * -2.1437327e-24 = -7.0616125e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011110111010000110100011011011;
		b = 32'b00111011100100011101111001110000;
		correct = 32'b11100010110010111111000010000010;
		#400 //-8.373438e+18 * 0.0044515654 = -1.8810097e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011000010011001010010000001111;
		b = 32'b00111100100110000000011100000110;
		correct = 32'b10011011001011000100110001001100;
		#400 //-2.644921e-24 * 0.018558037 = -1.425216e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110110111011010000001100000101;
		b = 32'b00111101110011111001000010011001;
		correct = 32'b01111000100100100010100011000001;
		#400 //2.4035852e+33 * 0.10135002 = 2.3715685e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110101111110110111110001010;
		b = 32'b11100110010000001111100000111111;
		correct = 32'b00001111111111011111011100000110;
		#400 //-5.7052284e-06 * -2.2781842e+23 = 2.5042876e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000010010010110100011011101;
		b = 32'b11000101010010100011110000011010;
		correct = 32'b00101010011111101111010010011010;
		#400 //-7.3272394e-10 * -3235.7563 = 2.2644595e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110000101101111100110101111110;
		b = 32'b11010101100100011111001101011011;
		correct = 32'b01011010101000010011001001010110;
		#400 //-4.5507345e+29 * -20059299000000.0 = 2.2686408e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001000100000010000000111000000;
		b = 32'b10010101100001111100010110000101;
		correct = 32'b00110010011100110011111010110111;
		#400 //-7.7643165e-34 * -5.4837697e-26 = 1.4158721e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000010100111111001110101010101;
		b = 32'b10001101001100101000100111000101;
		correct = 32'b11110100111001001101110110111000;
		#400 //79.80729 * -5.501632e-31 = -1.4506112e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111000100111000101101001110100;
		b = 32'b01101110010011011110110010000100;
		correct = 32'b00001001110000100101111111111111;
		#400 //7.455508e-05 * 1.5932589e+28 = 4.6794075e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010101110000000100000111011100;
		b = 32'b00101110010100000101000001001101;
		correct = 32'b00100110111011000100010010011101;
		#400 //7.765209e-26 * 4.7365046e-11 = 1.6394387e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101110110000100010001011110111;
		b = 32'b11001010100011100000011010000111;
		correct = 32'b01100011101011101111011100000110;
		#400 //-3.004118e+28 * -4653891.5 = 6.455067e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110110010111001001011011101011;
		b = 32'b01000101001100001011100011110011;
		correct = 32'b11110000100111111100010111011101;
		#400 //-1.1185218e+33 * 2827.5593 = -3.9557855e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100100101110111000111000110101;
		b = 32'b11100001010101100100011110111100;
		correct = 32'b10000010111000000001001001110010;
		#400 //8.133923e-17 * -2.4704826e+20 = -3.292443e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111110100001111000101110000111;
		b = 32'b10001111011001010101000110101001;
		correct = 32'b01101110100101110101000011001000;
		#400 //-0.26473638 * -1.1306299e-29 = 2.3414948e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010011010111001100011111001111;
		b = 32'b01111111011000010010010110100110;
		correct = 32'b00010011011110110000100011111010;
		#400 //948245040000.0 * 2.9927178e+38 = 3.168508e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010001101100010101001110001100;
		b = 32'b00111010110111000101111110111001;
		correct = 32'b10010110010011011111111001001000;
		#400 //-2.7977166e-28 * 0.0016813196 = -1.6640005e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010111111001100111100001010001;
		b = 32'b00000100110100110001010000100001;
		correct = 32'b01010010100010111100001001010100;
		#400 //1.4893774e-24 * 4.9624347e-36 = 300130370000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101010100001110011111011111011;
		b = 32'b01010010101100011010011010000101;
		correct = 32'b01010111010000101110010011010010;
		#400 //8.17512e+25 * 381501470000.0 = 214288030000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010111011111001011000101011110;
		b = 32'b00100010001011001110011000001111;
		correct = 32'b11110100101110110001001010110100;
		#400 //-277838720000000.0 * 2.3432139e-18 = -1.1857164e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110100111001010001010111101110;
		b = 32'b01001000011001001010110001011110;
		correct = 32'b01101100000000000011101100010111;
		#400 //1.4520029e+32 * 234161.47 = 6.200862e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111100100000011010001111000001;
		b = 32'b01101000100101101000111000011010;
		correct = 32'b01010011010111000110111110011011;
		#400 //5.385021e+36 * 5.68781e+24 = 946765230000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010110001000001000101011110010;
		b = 32'b01000001001100100111010101010101;
		correct = 32'b00010100011001100100110011001010;
		#400 //1.296854e-25 * 11.1536455 = 1.16271765e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101000101001111000010001101010;
		b = 32'b01001100010000000101110011111001;
		correct = 32'b10011011110111101110111101000100;
		#400 //-1.859815e-14 * 50426852.0 = -3.688144e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111000010011011101111100111111;
		b = 32'b01011011000000101001000010101001;
		correct = 32'b00011100110010011101001111010111;
		#400 //4.9083723e-05 * 3.6750802e+16 = 1.3355824e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010101000101000010100110001001;
		b = 32'b10001001000100100000101111000010;
		correct = 32'b01001011100000011101101011010101;
		#400 //-2.9921127e-26 * -1.757964e-33 = 17020330.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110101011110110111001001111100;
		b = 32'b01001000110111001001101101100110;
		correct = 32'b01101100000100011110010011011101;
		#400 //3.187472e+32 * 451803.2 = 7.055001e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100001100100001010000011110010;
		b = 32'b01011001101110101100101100111111;
		correct = 32'b01000111010001100011011001111001;
		#400 //3.3349106e+20 * 6572227000000000.0 = 50742.473
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000000001101011011100000101111;
		b = 32'b00110011010010011011011100010100;
		correct = 32'b00001100000010000101101000111110;
		#400 //4.933354e-39 * 4.6965468e-08 = 1.0504215e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100001111001001011000100101101;
		b = 32'b00100000011000010101101001011110;
		correct = 32'b01000001000000011110010110001000;
		#400 //1.5496779e-18 * 1.9088141e-19 = 8.118538
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001001001110001000111010111001;
		b = 32'b11111011001010010010110001001110;
		correct = 32'b10001101100010111010001111100100;
		#400 //755947.56 * -8.783968e+35 = -8.605992e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001100001000110001101101110101;
		b = 32'b11111011000011000001010101111011;
		correct = 32'b00010000100101010000100110001101;
		#400 //-42757588.0 * -7.273572e+35 = 5.878485e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010011101100110111001110011000;
		b = 32'b00010001010000011010001011100101;
		correct = 32'b11000001111011010011111100101110;
		#400 //-4.5299937e-27 * 1.5275211e-28 = -29.65585
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101100011001000011001001000101;
		b = 32'b01110110000101110010011000010111;
		correct = 32'b10110101110000010011111101100000;
		#400 //-1.1034899e+27 * 7.664154e+32 = -1.4398065e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011011101011111001101011001110;
		b = 32'b01001001010100010011011010001100;
		correct = 32'b01010001110101101110000000101110;
		#400 //9.885666e+16 * 856936.75 = 115360510000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101101011110110010110000001000;
		b = 32'b00111111000101111001000001001011;
		correct = 32'b11101101110101000001111101001001;
		#400 //-4.858373e+27 * 0.5920455 = -8.2060804e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010010010111001101000011101101;
		b = 32'b00110111001101111000111100000011;
		correct = 32'b11011010100110011111101100000110;
		#400 //-237099500000.0 * 1.09409475e-05 = -2.1670837e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101100000101111001100011001000;
		b = 32'b00011011101111001100010100110010;
		correct = 32'b11001111110011011001011001011011;
		#400 //-2.1543201e-12 * 3.1229426e-22 = -6898366000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110010001011011001101011010110;
		b = 32'b01100011010000110100010011001011;
		correct = 32'b00001110011000111001100100101100;
		#400 //1.0105131e-08 * 3.6020722e+21 = 2.805366e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101101110001100010000011111000;
		b = 32'b10011111000011000101001111011001;
		correct = 32'b01001110001101001011100100111000;
		#400 //-2.2524635e-11 * -2.971551e-20 = 758009340.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100000010000001110010101001;
		b = 32'b10110101101100100100001000011110;
		correct = 32'b11001101110000110111100100010000;
		#400 //544.4478 * -1.3281276e-06 = -409936400.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000000001110110110011110101100;
		b = 32'b00001000100101011111101101110000;
		correct = 32'b11110111000111111111000000011011;
		#400 //-2.9282026 * 9.026724e-34 = -3.2439262e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110001010100001010110010011000;
		b = 32'b00110010010010011100101100100011;
		correct = 32'b11111110100001000101110101010000;
		#400 //-1.03330456e+30 * 1.1745928e-08 = -8.79713e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001101011000100111101011100011;
		b = 32'b10111011101000100111110110011111;
		correct = 32'b11010001001100100110100000100011;
		#400 //237481520.0 * -0.004958823 = -47890706000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010101010010011010000101111011;
		b = 32'b00011000110010101111100011110101;
		correct = 32'b01111011111111100100111011001010;
		#400 //13855962000000.0 * 5.246716e-24 = 2.6408829e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010100010111100101110110111010;
		b = 32'b10011100101011110100011000101111;
		correct = 32'b10110111001000100110001111111010;
		#400 //1.122662e-26 * -1.1598671e-21 = -9.67923e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011000011110110000000101011001;
		b = 32'b00101010110011011010111110011110;
		correct = 32'b11101101000111000011001111011001;
		#400 //-1103932800000000.0 * 3.6537174e-13 = -3.0213963e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111111000110101100111010100110;
		b = 32'b00101101110111110100111111001100;
		correct = 32'b01010000101100010111011111000101;
		#400 //0.6047157 * 2.5387602e-11 = 23819332000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100100000011100111111011000000;
		b = 32'b11000000101110100000010000010100;
		correct = 32'b00100010110001000001101100000011;
		#400 //-3.0898703e-17 * -5.812998 = 5.3154506e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010011100111111110010111110010;
		b = 32'b10011000111100100001000101111010;
		correct = 32'b10111010001010010001100111010000;
		#400 //4.0363986e-27 * -6.257318e-24 = -0.0006450685
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001111111100100011010001001011;
		b = 32'b10100011010100110000001110010111;
		correct = 32'b00101100000100101110101101111011;
		#400 //-2.3883185e-29 * -1.1439093e-17 = 2.0878566e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001110100101110100110101010111;
		b = 32'b01011110011011101101001111100011;
		correct = 32'b00101111101000100010111001011110;
		#400 //1269214100.0 * 4.302337e+18 = 2.9500574e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011000001110111100000001000010;
		b = 32'b10100011110110100101100110011011;
		correct = 32'b10110011110111000001111111110100;
		#400 //2.4266249e-24 * -2.3673557e-17 = -1.02503606e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001110010011001110100110101110;
		b = 32'b10110000010110111100101101001001;
		correct = 32'b11011101011011101010101011011010;
		#400 //859466600.0 * -7.996062e-10 = -1.07486236e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001001100001101110101000001011;
		b = 32'b10100011110100100001111001010010;
		correct = 32'b10100101001001000101111111001001;
		#400 //3.247942e-33 * -2.2781087e-17 = -1.4257186e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000000010011111110001001110111;
		b = 32'b11101010101111000010010100101000;
		correct = 32'b10010101000011010110110111100101;
		#400 //3.2481973 * -1.1372676e+26 = -2.8561415e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100010110001001101100101100111;
		b = 32'b10011101100011001101010110101111;
		correct = 32'b11000100101100101110100011100101;
		#400 //5.335609e-18 * -3.7278635e-21 = -1431.278
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010010101100101110011101000010;
		b = 32'b01001001111011000100110010110111;
		correct = 32'b11001000010000011101000110001100;
		#400 //-384192020000.0 * 1935766.9 = -198470.19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110010001101001100101110011101;
		b = 32'b01000100010100111111001001001001;
		correct = 32'b11101101010110100101111111000110;
		#400 //-3.581021e+30 * 847.7857 = -4.2239697e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100111100100101010100001001101;
		b = 32'b10010111100010000001001001000011;
		correct = 32'b01001111100010011111010101001010;
		#400 //-4.0705612e-15 * -8.793404e-25 = 4629107700.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000010010100000111011000111111;
		b = 32'b10110101001111110001101101000000;
		correct = 32'b00001100100010111001111111011001;
		#400 //-1.5315362e-37 * -7.11927e-07 = 2.1512546e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100011111000101100011111011110;
		b = 32'b00100101000101001111011000001111;
		correct = 32'b01111110010000101101111010000000;
		#400 //8.366732e+21 * 1.2920322e-16 = 6.475638e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101001010111110000100111010011;
		b = 32'b11001000101001100100100011111111;
		correct = 32'b01100000001010111010111110111110;
		#400 //-1.6852303e+25 * -340551.97 = 4.9485262e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010010110111111101010101011111;
		b = 32'b00010110110011101011011000001000;
		correct = 32'b00111011100010101001101001000010;
		#400 //1.4125879e-27 * 3.3395973e-25 = 0.0042298147
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011000001010100000011000111011;
		b = 32'b00110011011010011110111000011100;
		correct = 32'b10100100001110100001000010101010;
		#400 //-2.197513e-24 * 5.44661e-08 = -4.0346436e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101001110010011110011100000111;
		b = 32'b00101011111000010010111011011011;
		correct = 32'b10111101011001011000100010001101;
		#400 //-8.96627e-14 * 1.6000217e-12 = -0.056038428
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101000110101010101111110110110;
		b = 32'b11001010000000011010101001001100;
		correct = 32'b11011110010100101010001000110101;
		#400 //8.061037e+24 * -2124435.0 = -3.794438e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011101100101010100101000000010;
		b = 32'b10111100101001100011101110110111;
		correct = 32'b01100000011001011110011111101001;
		#400 //-1.3446766e+18 * -0.020292146 = 6.6265864e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010111010100100111101000000100;
		b = 32'b01000111011000011001110000111100;
		correct = 32'b11001111011011101101001111101101;
		#400 //-231421500000000.0 * 57756.234 = -4006866200.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000011000111010010111010001110;
		b = 32'b01110111001111000100101100010111;
		correct = 32'b00001011010101011011001110010010;
		#400 //157.18185 * 3.8190422e+33 = 4.1157402e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101111100110010001000010111000;
		b = 32'b01100100001111101111110100101101;
		correct = 32'b00001010110011010010101011011110;
		#400 //2.7842417e-10 * 1.4092498e+22 = 1.9756907e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100001111100101101000110001101;
		b = 32'b00010001101010111010110101100010;
		correct = 32'b11001111101101010000101010111000;
		#400 //-1.6454025e-18 * 2.7085898e-28 = -6074757000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110011010100100101001010000001;
		b = 32'b11001001001010011001100101110111;
		correct = 32'b01101001100111101011101111111010;
		#400 //-1.6663448e+31 * -694679.44 = 2.3987247e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101010110011100010001001011010;
		b = 32'b10110110001011100000101100110100;
		correct = 32'b11110100000101111001100111001111;
		#400 //1.2460047e+26 * -2.5934542e-06 = -4.8044216e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010001110111000011101000001001;
		b = 32'b11110000011110010000001100000101;
		correct = 32'b10100000111000100110100000110111;
		#400 //118233310000.0 * -3.0826167e+29 = -3.8354853e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000001110001001101000000101110;
		b = 32'b00101100111111001111001010000001;
		correct = 32'b01010100010001110011000000111111;
		#400 //24.60165 * 7.189194e-12 = 3422031700000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001001001010000100010101110000;
		b = 32'b00010100110110000011010111100001;
		correct = 32'b01110011110001110011110100001011;
		#400 //689239.0 * 2.1831678e-26 = 3.1570592e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010011110101001001010111001101;
		b = 32'b11001011101011101010110100000011;
		correct = 32'b10000111100110111100011110001001;
		#400 //5.366404e-27 * -22895110.0 = -2.3439084e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100011100111111101100010111001;
		b = 32'b00001100100111100001010000100001;
		correct = 32'b11010110100000010110111001111010;
		#400 //-1.73306e-17 * 2.435587e-31 = -71155750000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010010001111000000100100011111;
		b = 32'b01000010010011100001101011010011;
		correct = 32'b10001111011010011000111001111010;
		#400 //-5.9333583e-28 * 51.526196 = -1.1515227e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010100111000000110100011100;
		b = 32'b10010000001100110000100011001100;
		correct = 32'b01101001110111110010001011110101;
		#400 //-0.0011905762 * -3.5308302e-29 = 3.3719442e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100010110100001000011000000111;
		b = 32'b00110010001100010000001010010110;
		correct = 32'b01110000000101101100100111000000;
		#400 //1.9232902e+21 * 1.0303344e-08 = 1.866666e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001001111000000111100010001010;
		b = 32'b00110011110111111001011000000110;
		correct = 32'b00010101100000001000000110101101;
		#400 //5.4039393e-33 * 1.0411536e-07 = 5.190338e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100101001100001111110100000101;
		b = 32'b00110001011010011101010111100101;
		correct = 32'b11110011010000011100001110110101;
		#400 //-5.2237743e+22 * 3.4027547e-09 = -1.5351604e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111101101001011100101100010;
		b = 32'b10011010000111010000100010000010;
		correct = 32'b11101101000100110100111110010001;
		#400 //92530.766 * -3.2473712e-23 = -2.8494054e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001100000111100000010110100011;
		b = 32'b01110101010110001000101000000100;
		correct = 32'b10010110001110101101000110101110;
		#400 //-41424524.0 * 2.7449595e+32 = -1.5091124e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000001011001101100000000000100;
		b = 32'b00101000001110011001001000111011;
		correct = 32'b10011000100111110010100110100100;
		#400 //-4.2382093e-38 * 1.0301272e-14 = -4.1142583e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110111011011001110101110111000;
		b = 32'b11000101000001101110111110101110;
		correct = 32'b10110001111000001011110111111100;
		#400 //1.4121579e-05 * -2158.98 = -6.5408567e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101101001111001011010011011111;
		b = 32'b11011010001010100100010001000011;
		correct = 32'b11010010100011011101110011000110;
		#400 //3.650115e+27 * -1.198145e+16 = -304647180000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010101010100111100100100010000;
		b = 32'b01101100100100000001111101100111;
		correct = 32'b10101000001111000001011111101101;
		#400 //-14553782000000.0 * 1.3938689e+27 = -1.04412845e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001011111000011110010100011000;
		b = 32'b01000001011001100010101110011101;
		correct = 32'b00001001111110110011111010100111;
		#400 //8.701155e-32 * 14.385648 = 6.048497e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100001010001111101001011011101;
		b = 32'b11110010111111111101011001000011;
		correct = 32'b10101101110001111111001101110111;
		#400 //2.3038102e+20 * -1.0134746e+31 = -2.27318e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111110101111101011010100001111;
		b = 32'b10110100110110000010110000011100;
		correct = 32'b01001001011000011101011111100000;
		#400 //-0.37247512 * -4.026523e-07 = 925054.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101111001100100100101110001100;
		b = 32'b11011100000001000111110011000101;
		correct = 32'b00010010101011000100000110010111;
		#400 //-1.6215845e-10 * -1.4916753e+17 = 1.0870895e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100001010100100100111010011010;
		b = 32'b00111001100010111011001001110000;
		correct = 32'b01100111010000001011001010011111;
		#400 //2.424675e+20 * 0.00026645092 = 9.0998934e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110011111001010101001000110100;
		b = 32'b01101110011010110001100110101100;
		correct = 32'b11000100111110011011010100000011;
		#400 //-3.633738e+31 * 1.8190003e+28 = -1997.6566
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100000111100000111111111011100;
		b = 32'b00100110110101111100000110111100;
		correct = 32'b11111001100011101010110111001001;
		#400 //-1.3863849e+20 * 1.4971134e-15 = -9.260387e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011000111011011100001010101111;
		b = 32'b10101001100101101011010011111000;
		correct = 32'b11101110110010011110111111110001;
		#400 //2091363300000000.0 * -6.692731e-14 = -3.124828e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111011111010010100100010011011;
		b = 32'b11000100011101011111000001010010;
		correct = 32'b10110110111100101101001111000000;
		#400 //0.007119251 * -983.755 = -7.236813e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100101010000101100001010100011;
		b = 32'b10110100110000101101110011100101;
		correct = 32'b10101111111111111101110110000001;
		#400 //1.6892763e-16 * -3.6296038e-07 = -4.6541618e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110111110101110001110101000111;
		b = 32'b00001010010100111011101111101100;
		correct = 32'b01101101000000100000101100100011;
		#400 //2.564363e-05 * 1.0194625e-32 = 2.5154072e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100101000011011010100000011000;
		b = 32'b11011110101010000111100110100111;
		correct = 32'b01000101110101110011111110110101;
		#400 //-4.1809654e+22 * -6.069959e+18 = 6887.9634
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101011111100101110000010100011;
		b = 32'b00111011010110001000101100011111;
		correct = 32'b10110000000011111001000011110010;
		#400 //-1.7257483e-12 * 0.0033041907 = -5.2229077e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010001110101110111001101011;
		b = 32'b10101000111011100111010010110000;
		correct = 32'b01010000110010001010111101000100;
		#400 //-0.0007130864 * -2.6473913e-14 = 26935435000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111101100010011111110101101010;
		b = 32'b11001110001010000110111000001010;
		correct = 32'b00101110110100011011101111010100;
		#400 //-0.06737788 * -706445950.0 = 9.5375846e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010110001111101011111011001111;
		b = 32'b00100100101001111111010011000000;
		correct = 32'b01110001000100010101111000101001;
		#400 //52431680000000.0 * 7.283933e-17 = 7.1982655e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110011000011111100011111001000;
		b = 32'b01011010101101101101100101010110;
		correct = 32'b01010111110010010100110100110011;
		#400 //1.1391457e+31 * 2.5733705e+16 = 442666800000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110010000110010011011001010110;
		b = 32'b10010111010001001101001010010110;
		correct = 32'b11011010010001110100011100010001;
		#400 //8.918127e-09 * -6.3596812e-25 = -1.4022915e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001101010101001001101010000110;
		b = 32'b10000010100110000100100011110111;
		correct = 32'b11001010001100101011001100010101;
		#400 //6.5513545e-31 * -2.2376272e-37 = -2927813.2
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100000101111111010011101000110;
		b = 32'b11010100100111100010010100011100;
		correct = 32'b10001011100110110001111100000111;
		#400 //3.246735e-19 * -5433819400000.0 = -5.9750513e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110010100001100001010111111;
		b = 32'b00101111110101100010001100010111;
		correct = 32'b01001101111110011001001010010110;
		#400 //0.2038679 * 3.8951306e-10 = 523391680.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010110110111011101100101010010;
		b = 32'b00010111001001111001000101101001;
		correct = 32'b11111111001010010111011010101000;
		#400 //-121962730000000.0 * 5.4144144e-25 = -2.2525563e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010001010101111010100001011101;
		b = 32'b10111011111111000011001100111010;
		correct = 32'b01010100110110101110100000110000;
		#400 //-57890165000.0 * -0.0076965364 = 7521586600000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001100010011011111010010101100;
		b = 32'b01000100110110101101111010100100;
		correct = 32'b11000110111100001110010100110000;
		#400 //-53990064.0 * 1750.9575 = -30834.594
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100110000100010110000100100000;
		b = 32'b00001101100110100100111011010101;
		correct = 32'b11010111111100010010111111110111;
		#400 //-5.043861e-16 * 9.509961e-31 = -530376620000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001101001101101000010011101011;
		b = 32'b00100110100100010110100000111000;
		correct = 32'b01100110001000001010101101011000;
		#400 //191385260.0 * 1.0089645e-15 = 1.8968484e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000011101000110111101010011011;
		b = 32'b00110111000110000111100001000000;
		correct = 32'b11001100000010010011111000001010;
		#400 //-326.95786 * 9.087904e-06 = -35977256.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111010011110011100000110111000;
		b = 32'b11101010001010011011110000111100;
		correct = 32'b11001111101111000101100001101011;
		#400 //3.2420275e+35 * -5.1299344e+25 = -6319822300.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101101001100100101110110000100;
		b = 32'b01011100000110111000001000011010;
		correct = 32'b10010000100100101101000001011000;
		#400 //-1.0138893e-11 * 1.7508668e+17 = -5.790785e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100110110100010110011110111100;
		b = 32'b10110001110101100000111100110000;
		correct = 32'b10110100011110100110111100011011;
		#400 //1.4530406e-15 * -6.2299463e-09 = -2.3323484e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100100001110101101110100011000;
		b = 32'b11100001100010100110011111001011;
		correct = 32'b11000010001011001101000010101001;
		#400 //1.3788104e+22 * -3.1914122e+20 = -43.20377
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011111100100111110110101001001;
		b = 32'b00110101000000101001000100000111;
		correct = 32'b11101010000100010000010011100110;
		#400 //-2.1318512e+19 * 4.8639816e-07 = -4.3829344e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110010011101101011100001000000;
		b = 32'b01101111101001101000111010101011;
		correct = 32'b01000010001111011001101011101101;
		#400 //4.8867876e+30 * 1.0309397e+29 = 47.401295
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000001101110010101101000110001;
		b = 32'b01101010101000000100101110111011;
		correct = 32'b00010110100101000000001000011001;
		#400 //23.169039 * 9.689288e+25 = 2.3912013e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110001110111101011001010010100;
		b = 32'b01000110111101111011001110011011;
		correct = 32'b00101010011001100010100010000111;
		#400 //6.4813523e-09 * 31705.803 = 2.0442164e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100101101100000011010000101010;
		b = 32'b01011111110010100101111011110101;
		correct = 32'b10000101010111101110011000000000;
		#400 //-3.056648e-16 * 2.9164724e+19 = -1.0480634e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100110001001101101011110010000;
		b = 32'b10100111100100111001110110101010;
		correct = 32'b00111110000100001010101111011011;
		#400 //-5.788496e-16 * -4.0971636e-15 = 0.14128058
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001001000111011000010010001100;
		b = 32'b10010110111100110111100111011101;
		correct = 32'b01110001101001011001111011000101;
		#400 //-645192.75 * -3.9335674e-25 = 1.640223e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100000001111101110011001000110;
		b = 32'b11110101110001100101010001110011;
		correct = 32'b00101001111101100110100010110110;
		#400 //-5.5023036e+19 * -5.02826e+32 = 1.0942759e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011110001110000010100111000111;
		b = 32'b10110110010101111010001100000111;
		correct = 32'b11100111010110101010001010010101;
		#400 //3.3175891e+18 * -3.213239e-06 = -1.032475e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010000010111101001000001000101;
		b = 32'b00011101100110111110001000100111;
		correct = 32'b00110010001101101100000010111010;
		#400 //4.389292e-29 * 4.1261994e-21 = 1.0637615e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111001001111000101000111111000;
		b = 32'b01001000111111010101001011011101;
		correct = 32'b10101111101111100100111101001100;
		#400 //-0.00017959613 * 518806.9 = -3.4617142e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111100110100110110001011010010;
		b = 32'b11001101111111111010101110100000;
		correct = 32'b11101110010100111010100010010101;
		#400 //8.7806316e+36 * -536179700.0 = -1.6376285e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011000010111111010001100100000;
		b = 32'b10011011101000011100010000000011;
		correct = 32'b11111100001100001111010011111100;
		#400 //983566840000000.0 * -2.6761885e-22 = -3.6752525e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110011010001001001101000011110;
		b = 32'b11100001110101011000011111100011;
		correct = 32'b00010000111010111011010001001001;
		#400 //-4.5774975e-08 * -4.9236852e+20 = 9.296893e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100110111100011001110110110111;
		b = 32'b10111111100111011101001000011001;
		correct = 32'b00100110110000111111011001000101;
		#400 //-1.6765483e-15 * -1.2329742 = 1.3597595e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001000111110000010110000011010;
		b = 32'b11111010011101100111111101100111;
		correct = 32'b10001110000000001101111010011101;
		#400 //508256.8 * -3.1997226e+35 = -1.5884403e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100010100000000101010011111001;
		b = 32'b11101001101101100000111000001110;
		correct = 32'b10111000001101000111010011010111;
		#400 //1.1836531e+21 * -2.7511359e+25 = -4.302416e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110001101011001011100111110;
		b = 32'b01111011101010100100100000100110;
		correct = 32'b00000010000010001000000000111010;
		#400 //0.17733476 * 1.7683076e+36 = 1.0028501e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011010001010100111111100011110;
		b = 32'b11010010110110110100011011101001;
		correct = 32'b01000110110001110000110011010110;
		#400 //-1.1997628e+16 * -470893760000.0 = 25478.418
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110111101011111110110001100101;
		b = 32'b11101010010001000000111011011111;
		correct = 32'b10001100111001011011010110011110;
		#400 //2.0971705e-05 * -5.925492e+25 = -3.5392343e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111011110100011101100101000101;
		b = 32'b01101111110001110010001010011101;
		correct = 32'b11001011100001101110001011101100;
		#400 //-2.1791936e+36 * 1.2325872e+29 = -17679832.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001111100100011100111111000001;
		b = 32'b10110100101001010110001100101110;
		correct = 32'b11011010011000011011001011101001;
		#400 //4892623400.0 * -3.0805808e-07 = -1.5882146e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111110100010101101010101000111;
		b = 32'b01111101011111111000101000010001;
		correct = 32'b11000000100010110001010101011010;
		#400 //-9.227043e+37 * 2.1229376e+37 = -4.3463564
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001010101001100110000010110010;
		b = 32'b10010110001010110001001010110000;
		correct = 32'b11110011111110001111100101001011;
		#400 //5451865.0 * -1.3819167e-25 = -3.9451473e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011000001001111000100111101000;
		b = 32'b11001101001011100110111110111000;
		correct = 32'b11001010011101011110000010000110;
		#400 //736843000000000.0 * -182909820.0 = -4028449.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110010101111111101111110101110;
		b = 32'b01010110100001011110000010100100;
		correct = 32'b11011011101101110111001100111001;
		#400 //-7.600902e+30 * 73599935000000.0 = -1.0327322e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110010001010100001110001110000;
		b = 32'b01110110000110010011010010010000;
		correct = 32'b10111011100011100001111111011010;
		#400 //-3.3693972e+30 * 7.768433e+32 = -0.004337293
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110010100001001101010110100001;
		b = 32'b00000001000101000110000101010110;
		correct = 32'b01110000111001010010110111010010;
		#400 //1.546397e-08 * 2.7253142e-38 = 5.674197e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010100111110100011011110110100;
		b = 32'b10100001001111011001110111000111;
		correct = 32'b00110011001010001110100010100011;
		#400 //-2.526552e-26 * -6.4244507e-19 = 3.932713e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000100001001100110000000101011;
		b = 32'b11001011001100101101111101111100;
		correct = 32'b00111000011011100001110100110001;
		#400 //-665.5026 * -11722620.0 = 5.677081e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110011011101010110001110100101;
		b = 32'b01000100001100111000000001111110;
		correct = 32'b11101110101011101111101110110100;
		#400 //-1.9441738e+31 * 718.0077 = -2.707734e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111000001000000011001011101101;
		b = 32'b10111101011001100111011011110011;
		correct = 32'b00111010001100011111001011101010;
		#400 //-3.81944e-05 * -0.056265783 = 0.0006788211
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010100110111001101001100011110;
		b = 32'b10100111001000011011110100001100;
		correct = 32'b10101101001011101100001011001010;
		#400 //2.2297594e-26 * -2.244572e-15 = -9.934007e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001010010111010111010100010001;
		b = 32'b00011111001101111001100010100001;
		correct = 32'b01101010100110100110010101100101;
		#400 //3628356.2 * 3.887801e-20 = 9.33267e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010111111110010101011111001101;
		b = 32'b11111010110011010100010100011010;
		correct = 32'b10011100100110110111101110001011;
		#400 //548311000000000.0 * -5.329112e+35 = -1.0288975e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001100101101101100101100000010;
		b = 32'b00110111000101011010010111010110;
		correct = 32'b10010101000111000101100110111001;
		#400 //-2.816372e-31 * 8.919704e-06 = -3.1574728e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111110111010011000100000111;
		b = 32'b01101111101011101111001010000111;
		correct = 32'b00010111101000011101010110011111;
		#400 //113250.055 * 1.0828718e+29 = 1.0458307e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010001111111111010010001101001;
		b = 32'b00101100101000001100111010100000;
		correct = 32'b00100100110010110111110010111110;
		#400 //4.0333232e-28 * 4.5704135e-12 = 8.824854e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011111011100010101111011001000;
		b = 32'b00100100001010010010000110100101;
		correct = 32'b01111010101101101010101111000001;
		#400 //1.7392559e+19 * 3.667453e-17 = 4.742408e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011001101000001000011001011000;
		b = 32'b10101110111011100000001000111000;
		correct = 32'b00101010001011001010100010110110;
		#400 //-1.6597873e-23 * -1.0823381e-10 = 1.5335202e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100001111111111111010111000001;
		b = 32'b11010011000110010000001010010110;
		correct = 32'b01001110010101100001111101010000;
		#400 //-5.9020352e+20 * -657173400000.0 = 898094100.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001110111111100110001001001000;
		b = 32'b00100001001110101001010101010100;
		correct = 32'b10101101001011101000001100111010;
		#400 //-6.2710476e-30 * 6.3216885e-19 = -9.919893e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001101100110011101011010010110;
		b = 32'b01100011100001000101111010110111;
		correct = 32'b00101001100101001100001001101111;
		#400 //322622140.0 * 4.8835903e+21 = 6.606249e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000100010111011111010011100101;
		b = 32'b00001010010100011000001101011100;
		correct = 32'b00111001100001111001101000101100;
		#400 //2.6090875e-36 * 1.008769e-32 = 0.00025864074
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000000000100100011011001001101;
		b = 32'b00111010001111001110000100001011;
		correct = 32'b01000101010001100010101110110100;
		#400 //2.2845643 * 0.0007205165 = 3170.7314
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011100001110000101011101000000;
		b = 32'b01000111011111100111101011110110;
		correct = 32'b11010100001110010111000100010000;
		#400 //-2.0754931e+17 * 65146.96 = -3185863300000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010101110111011100000010100010;
		b = 32'b00110001110001100111010101111101;
		correct = 32'b11100011100011110000011000001100;
		#400 //-30477428000000.0 * 5.7759153e-09 = -5.27664e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000011001111000111000111010001;
		b = 32'b01011100111010111010111100010111;
		correct = 32'b10100101110011001011000001001000;
		#400 //-188.4446 * 5.3071306e+17 = -3.5507812e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010100111101110110111110000100;
		b = 32'b00110000110000001111101000100011;
		correct = 32'b10100011101001000001111100110001;
		#400 //-2.4984612e-26 * 1.4040932e-09 = -1.7794126e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100001000110101101111101100100;
		b = 32'b11010110101001111111101011001101;
		correct = 32'b11001001111011000000011001100000;
		#400 //1.7855597e+20 * -92347810000000.0 = -1933516.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110001100110100001000110000011;
		b = 32'b00011111111110011000111100001011;
		correct = 32'b11010001000111100000101110000100;
		#400 //-4.4839807e-09 * 1.05692247e-19 = -42424877000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100001001001001001111111110101;
		b = 32'b01001101001000101110000100010001;
		correct = 32'b00010011100000010101111100110001;
		#400 //5.5777063e-19 * 170791180.0 = 3.2658044e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100000011001010000001110000110;
		b = 32'b11010100101111111101100001010010;
		correct = 32'b10001011000110001100110010011000;
		#400 //1.939822e-19 * -6591744000000.0 = -2.9428054e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010001110100001000010010111000;
		b = 32'b00100001010100101100110110011111;
		correct = 32'b10101111111111010011100110110001;
		#400 //-3.2898408e-28 * 7.1422905e-19 = -4.6061424e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101010101101011110000101011100;
		b = 32'b00000111010110011110010110111011;
		correct = 32'b11100010110101011010111101001111;
		#400 //-3.2308433e-13 * 1.6392777e-34 = -1.9708944e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110011111000010110011110000000;
		b = 32'b10110000101100010000100010000001;
		correct = 32'b11000010101000101111100101000001;
		#400 //1.04962055e-07 * -1.2880862e-09 = -81.486824
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001010000011010110001001001100;
		b = 32'b00111010110101111001010101100111;
		correct = 32'b11001110101001111110001111001101;
		#400 //-2316435.0 * 0.0016447724 = -1408362100.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110100111001000010100101011011;
		b = 32'b10101011111000111010000100100011;
		correct = 32'b11001000100000000100110010011001;
		#400 //4.24984e-07 * -1.6174045e-12 = -262756.78
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110010111100110011100010010011;
		b = 32'b01101000110110100000011001010100;
		correct = 32'b11001001100011101100101011011111;
		#400 //-9.634976e+30 * 8.236741e+24 = -1169755.9
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000011111110011111010100100100;
		b = 32'b01101111101001011111110000001111;
		correct = 32'b10010011110000001100000110011010;
		#400 //-499.91516 * 1.0273949e+29 = -4.865852e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110111110000011101110011101;
		b = 32'b10110110101000100101100100010100;
		correct = 32'b00111111110000111011011011011000;
		#400 //-7.397916e-06 * -4.8383463e-06 = 1.5290174
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100110001000100011001100001111;
		b = 32'b10011010001100100111100100101111;
		correct = 32'b01001011011010001010100000101001;
		#400 //-5.627424e-16 * -3.690743e-23 = 15247401.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100101011100101101101010011101;
		b = 32'b00011110100001100100001110000100;
		correct = 32'b11000110011001111000011000110100;
		#400 //-2.1064223e-16 * 1.4215726e-20 = -14817.551
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111110011010100101010100111010;
		b = 32'b11100110110010111011100101011101;
		correct = 32'b11010111000100110011101101000111;
		#400 //7.787047e+37 * -4.8102987e+23 = -161882800000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011101010111101110111101110100;
		b = 32'b11011000000000110001110010101010;
		correct = 32'b11000100110110011010010011011010;
		#400 //1.0040116e+18 * -576636540000000.0 = -1741.1516
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010110010011100101011011100101;
		b = 32'b11110101000110101001011100100010;
		correct = 32'b00100000101010101101100100010100;
		#400 //-56718150000000.0 * -1.9596657e+32 = 2.894277e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110111010010101110011111011;
		b = 32'b01100110011101100001100111110010;
		correct = 32'b10001111111100101011111111100000;
		#400 //-6.9547655e-06 * 2.9054519e+23 = -2.393695e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000011100011100101100101000001;
		b = 32'b10100111110000001111001111110001;
		correct = 32'b10011011001111001101110001100011;
		#400 //8.366502e-37 * -5.3555187e-15 = -1.5622206e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111101101001001100110011000111;
		b = 32'b11001001011110000010110011001001;
		correct = 32'b11110011101010011111111100000010;
		#400 //2.7382082e+37 * -1016524.56 = -2.693696e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110100110110010001010010101110;
		b = 32'b10001111100110010101101100100101;
		correct = 32'b01100100101101010011000000111101;
		#400 //-4.0434446e-07 * -1.5122072e-29 = 2.6738693e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101010011010100101110101101101;
		b = 32'b01100111111101110011111010000110;
		correct = 32'b01000001111100101010101000100100;
		#400 //7.083246e+25 * 2.3351558e+24 = 30.333076
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111001000110101110011000010011;
		b = 32'b00110100101100100001000101110110;
		correct = 32'b01000011110111101011000010111100;
		#400 //0.00014772294 * 3.3167788e-07 = 445.38074
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000000001100100011000100100100;
		b = 32'b10111101010001011000111011011011;
		correct = 32'b00000010000000100001010001100101;
		#400 //-4.609403e-39 * -0.04823194 = 9.556745e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010010011111001011111010000100;
		b = 32'b11100110100001100010001110110100;
		correct = 32'b10101011011100010010110100100001;
		#400 //271382020000.0 * -3.1672786e+23 = -8.568303e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010011100011001110010011011;
		b = 32'b00010000110100010000101100001110;
		correct = 32'b11101001000100111111000100110010;
		#400 //-0.00092167564 * 8.2453e-29 = -1.1178194e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100100100110100101011011001000;
		b = 32'b11100000110000000001010111010100;
		correct = 32'b01000011010011011011000110101000;
		#400 //-2.2776415e+22 * -1.1072962e+20 = 205.69397
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110010000110111101110010101010;
		b = 32'b01010011011101010110011111010110;
		correct = 32'b01011110001000101001011100110111;
		#400 //3.0871644e+30 * 1054009070000.0 = 2.9289734e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001000111000000110101110000111;
		b = 32'b10000010101110110110000111110111;
		correct = 32'b11000101100110010100110011001101;
		#400 //1.3506789e-33 * -2.753341e-37 = -4905.6
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010101001011011011100010000000;
		b = 32'b00001011000100011111101010100110;
		correct = 32'b01001001100110000101001100101100;
		#400 //3.5082617e-26 * 2.811455e-32 = 1247845.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110011101110000001000001001000;
		b = 32'b01001011110110111000110001000001;
		correct = 32'b00100111010101101001111111001010;
		#400 //8.571129e-08 * 28776578.0 = 2.9785088e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111101001001101011101011000101;
		b = 32'b11101110001100101010110100101001;
		correct = 32'b01001110011011101110001000010001;
		#400 //-1.3851351e+37 * -1.3824417e+28 = 1001948200.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011101000101100011010000001110;
		b = 32'b10000001000010110110100001111110;
		correct = 32'b01011011100010011110100101101010;
		#400 //-1.9879246e-21 * -2.5605237e-38 = 7.763743e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010001011011111111101000011110;
		b = 32'b11001000000000101101101101110101;
		correct = 32'b01001000111010101011110010110110;
		#400 //-64418340000.0 * -133997.83 = 480741.7
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000101010001100000000110010011;
		b = 32'b01010011100011001001010110110100;
		correct = 32'b10110001001101000100011111111010;
		#400 //-3168.0984 * 1207614000000.0 = -2.6234361e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100011100111111101011101010000;
		b = 32'b11010111011110001010010101010000;
		correct = 32'b11001011101001001001000110010111;
		#400 //5.8970944e+21 * -273388900000000.0 = -21570350.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110000101001111001001001000000;
		b = 32'b11110110010110001001110110111110;
		correct = 32'b00111001110001100000100110111111;
		#400 //-4.148864e+29 * -1.0983745e+33 = 0.00037772764
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000000000011011001010011001000;
		b = 32'b11001101011001101001011101111100;
		correct = 32'b10110010000111010010111001111110;
		#400 //2.212206 * -241792960.0 = -9.149174e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111001100000010111000100111;
		b = 32'b00101100001111011000100010000111;
		correct = 32'b01011010011011011111011011011001;
		#400 //45102.152 * 2.6934303e-12 = 1.6745245e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101000011101110011111011001001;
		b = 32'b10100000110000101110011011111101;
		correct = 32'b01000111001000100110000000101100;
		#400 //-1.3724869e-14 * -3.3017734e-19 = 41568.17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110101000111011010000010100000;
		b = 32'b10100101010111001100010011001111;
		correct = 32'b11001111001101101100100001000101;
		#400 //5.87208e-07 * -1.914864e-16 = -3066578200.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111100110010110101011000110110;
		b = 32'b01001010010110011111010010101101;
		correct = 32'b11110001111011101101010001001001;
		#400 //-8.4462786e+36 * 3570987.2 = -2.3652502e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011000101111011011101000011000;
		b = 32'b11001100101000111110101100101110;
		correct = 32'b01001011100101000010011100101101;
		#400 //-1668855700000000.0 * -85940590.0 = 19418714.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001011110110000111100001100110;
		b = 32'b10000011011100100100001100111011;
		correct = 32'b01000111111001001011111011000010;
		#400 //-8.338133e-32 * -7.1194585e-37 = 117117.516
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101101111100001000010001011000;
		b = 32'b11100110011011101010101110111001;
		correct = 32'b10000111000000001111110101111000;
		#400 //2.7343613e-11 * -2.8177274e+23 = -9.704137e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100111110001010011001010011010;
		b = 32'b11110101010110101111100101000001;
		correct = 32'b00110001111001101000101010111010;
		#400 //-1.8624793e+24 * -2.7758208e+32 = 6.7096524e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000100000100001010101000010100;
		b = 32'b00110110010101101011001110001000;
		correct = 32'b00001101001011000111110110111110;
		#400 //1.7005215e-36 * 3.1992986e-06 = 5.315295e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010111110110011100001111100010;
		b = 32'b11101010100011011111101010000110;
		correct = 32'b00101100110001000101001100101111;
		#400 //-478870670000000.0 * -8.58208e+25 = 5.5798903e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100010111011001001001101111100;
		b = 32'b00111010111000110011000011100000;
		correct = 32'b10100111100001010100100110100011;
		#400 //-6.4124083e-18 * 0.0017333291 = -3.6994753e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100101101000011010011011000110;
		b = 32'b11011001000001011101010010010011;
		correct = 32'b01001100000110101001101111101011;
		#400 //-9.542218e+22 * -2354368700000000.0 = 40529836.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001101101001000111011011010110;
		b = 32'b01111000001011110110100110110110;
		correct = 32'b00010100111100000000010101110010;
		#400 //344906430.0 * 1.4231188e+34 = 2.4235955e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001010011010011001111111000011;
		b = 32'b10001110010001100110111110001001;
		correct = 32'b11111011100101101011001010110111;
		#400 //3827696.8 * -2.4459086e-30 = -1.5649386e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010011010100110010010000100010;
		b = 32'b10010111101111011001001001000010;
		correct = 32'b11111011000011101001000001101001;
		#400 //906844300000.0 * -1.2250759e-24 = -7.4023514e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100001101111010111000010101110;
		b = 32'b01001000110000111011000001110011;
		correct = 32'b01011000011101111101001100110000;
		#400 //4.3681926e+20 * 400771.6 = 1089945660000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110010101000100000001010001001;
		b = 32'b10110110011011101010111001010110;
		correct = 32'b01111011101011011100001111111011;
		#400 //-6.4178735e+30 * -3.556624e-06 = 1.8044846e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000000111011000110110011101010;
		b = 32'b10111111011111111001111101101101;
		correct = 32'b10000000111011001100011000111100;
		#400 //2.1712248e-38 * -0.9985264 = -2.174429e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001111100110011101000010101000;
		b = 32'b10011101111001000101100101011111;
		correct = 32'b00110001001011000111000011001011;
		#400 //-1.5167336e-29 * -6.0443505e-21 = 2.509341e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000011110000011100100100111010;
		b = 32'b00011000010010000101010001011000;
		correct = 32'b01101010111101111010001101100000;
		#400 //387.57208 * 2.5891977e-24 = 1.496881e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100101010000010011011001011110;
		b = 32'b01100011111111001001011111110110;
		correct = 32'b11000000110000111101000101100111;
		#400 //-5.7026227e+22 * 9.319059e+21 = -6.119312
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101100111010101011100001101101;
		b = 32'b11001100011010001100101101010000;
		correct = 32'b01100000000000010000111100100010;
		#400 //-2.2700765e+27 * -61025600.0 = 3.7198757e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000100101110001010000111101110;
		b = 32'b10101011000000010010011011001110;
		correct = 32'b01011001001101101111110001111100;
		#400 //-1477.0603 * -4.588386e-13 = 3219128500000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101011001011101000101000000001;
		b = 32'b01101101010101001111101001101011;
		correct = 32'b10111101010100011100101111010000;
		#400 //-2.110048e+26 * 4.1195974e+27 = -0.05121976
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001110111001110010100000000100;
		b = 32'b10011000000100100000101001001001;
		correct = 32'b11110110010010101001101000010010;
		#400 //1939079700.0 * -1.887525e-24 = -1.0273134e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111010100110111110111010100101;
		b = 32'b01101000110010011010010110001000;
		correct = 32'b00010001010001011111011010100000;
		#400 //0.0011896683 * 7.6179934e+24 = 1.5616557e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010010000000000111010101100100;
		b = 32'b10111100110011011011110100100110;
		correct = 32'b00010100100111111101011100100111;
		#400 //-4.0534373e-28 * -0.025114607 = 1.613976e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011111000010100011011111100101;
		b = 32'b00001001101011001011101000111101;
		correct = 32'b11010100110011001101101010010111;
		#400 //-2.926887e-20 * 4.158263e-33 = -7038725000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001001011011010111100100100100;
		b = 32'b01110011111110101101111001101010;
		correct = 32'b00010100111100100101010010010110;
		#400 //972690.25 * 3.975175e+31 = 2.4469119e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000010101010000101101000100101;
		b = 32'b10011100100110010111000001101000;
		correct = 32'b00100101100011000111000011001001;
		#400 //-2.4737122e-37 * -1.0153747e-21 = 2.4362555e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111001011100110111110000010111;
		b = 32'b11010010011101000101011000100110;
		correct = 32'b11100110011111110001101110001000;
		#400 //7.901531e+34 * -262354340000.0 = -3.0117783e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010001010011001111001111011001;
		b = 32'b10110000000001111001101111100011;
		correct = 32'b00100000110000010111001111101001;
		#400 //-1.6167904e-28 * -4.933424e-10 = 3.2772175e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110010111000100110100010010110;
		b = 32'b11001101111011010100000001001100;
		correct = 32'b01100100011101000100110011110000;
		#400 //-8.968966e+30 * -497551740.0 = 1.8026198e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010000010011001101111010011010;
		b = 32'b10010111100101011000001100011010;
		correct = 32'b00111000001011110110010001111010;
		#400 //-4.0403392e-29 * -9.661994e-25 = 4.1816827e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000000111100011111011110100101;
		b = 32'b10110101100100101110011001001001;
		correct = 32'b01001010110100101101011000110100;
		#400 //-7.56148 * -1.094487e-06 = 6908698.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110001010010001010101101100100;
		b = 32'b01110111111011101000011010100010;
		correct = 32'b10111000110101110101111011001010;
		#400 //-9.936672e+29 * 9.6757604e+33 = -0.00010269655
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110100011010000010011111011111;
		b = 32'b00011000000011010100001000101101;
		correct = 32'b01011011110100100101110110011011;
		#400 //2.1621189e-07 * 1.8257233e-24 = 1.1842533e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001000100000101001000000111101;
		b = 32'b00110100110010111110111010010010;
		correct = 32'b00010011001000111110011000100101;
		#400 //7.858001e-34 * 3.798528e-07 = 2.0686962e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011110111011000111001001110011;
		b = 32'b10110010011011101111001110000100;
		correct = 32'b10101011111111010101000100110010;
		#400 //2.5034807e-20 * -1.3908792e-08 = -1.7999267e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010011001011111100010111110011;
		b = 32'b00111010000110100111011110110100;
		correct = 32'b01011000100100011010011110101101;
		#400 //754940300000.0 * 0.0005892471 = 1281194800000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111100011001011000100000100000;
		b = 32'b10100011001000011010010110100101;
		correct = 32'b11011000101101011100000100100000;
		#400 //0.0140095055 * -8.762904e-18 = -1598728600000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000011100001011000000010010111;
		b = 32'b00010001101111000111000001110101;
		correct = 32'b01110001001101010101110111011001;
		#400 //267.0046 * 2.9730477e-28 = 8.980839e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010010100110010000100000101111;
		b = 32'b00011101011011110100101100001101;
		correct = 32'b11110100101000111011011101011101;
		#400 //-328633650000.0 * 3.1670187e-21 = -1.0376751e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100001101011111011011110111;
		b = 32'b01001011000011000101001010000110;
		correct = 32'b00111000101001011111110001001100;
		#400 //727.8588 * 9196166.0 = 7.914807e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100100011111010110001111000001;
		b = 32'b11000001110000110011110001111101;
		correct = 32'b00100010001001100010000001010100;
		#400 //-5.4945125e-17 * -24.404535 = 2.251431e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010000110100001110010010000011;
		b = 32'b01000111001110000001000010101111;
		correct = 32'b00001001000100010100001111100001;
		#400 //8.239361e-29 * 47120.684 = 1.7485657e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001110111101100110101110000001;
		b = 32'b10000001101110010000000010101000;
		correct = 32'b11001100101010100111111001011100;
		#400 //6.0747205e-30 * -6.795921e-38 = -89387740.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010010011110001100011011010110;
		b = 32'b10010010011110101011101000011011;
		correct = 32'b10111111011111100000001000111011;
		#400 //7.8500086e-28 * -7.9115483e-28 = -0.99222153
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010011011010010111010011001000;
		b = 32'b11001011100101100000001101000101;
		correct = 32'b01000111010001110011001011110000;
		#400 //-1002686640000.0 * -19662474.0 = 50994.938
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010101110000100011010101010111;
		b = 32'b11101110011110101101110110000111;
		correct = 32'b00100110110001100010111011110010;
		#400 //-26691794000000.0 * -1.9409766e+28 = 1.3751734e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110111010110110011001101001001;
		b = 32'b01110101111100001101001000011111;
		correct = 32'b00000000111010010000010001001100;
		#400 //1.3065358e-05 * 6.1055323e+32 = 2.1399212e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010010111100000110111010100001;
		b = 32'b10111000100010100001000011011100;
		correct = 32'b01011001110111101110011100110101;
		#400 //-516324100000.0 * -6.583493e-05 = 7842707500000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101111010110000000000001000001;
		b = 32'b10010001001111101000101101010010;
		correct = 32'b11011101100100010001100111010001;
		#400 //1.9645176e-10 * -1.5031289e-28 = -1.3069522e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101100001100011111001000110111;
		b = 32'b11001011001111110011110111001100;
		correct = 32'b00100000011011100011001111100100;
		#400 //-2.528767e-12 * -12533196.0 = 2.0176553e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111101100010100000001110110101;
		b = 32'b00101101000011000101101111100111;
		correct = 32'b11001111111110111011100101001111;
		#400 //-0.06738988 * 7.978485e-12 = -8446451000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111101011010001111000010100000;
		b = 32'b11101101010011010010011111011101;
		correct = 32'b00001111100100010101010111000101;
		#400 //-0.056870103 * -3.9682887e+27 = 1.4331141e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100100111100000110110011100001;
		b = 32'b10110011100011110011011110101110;
		correct = 32'b00110000110101101110000100001001;
		#400 //-1.04267857e-16 * -6.6690845e-08 = 1.5634508e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100011100100100000000101001100;
		b = 32'b11111011101000111000011110011010;
		correct = 32'b10100111011001001001000011011001;
		#400 //5.386636e+21 * -1.6981894e+36 = -3.1719878e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111111110111101011001100111101;
		b = 32'b10100011000011110000000101011011;
		correct = 32'b01011100010001110101010100100110;
		#400 //-1.7398449 * -7.7523326e-18 = 2.2442857e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100001000011100101010010010110;
		b = 32'b00110111011001000011110000001111;
		correct = 32'b10101001000111111010010100110100;
		#400 //-4.822342e-19 * 1.36038425e-05 = -3.5448383e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000100011000011000010111011100;
		b = 32'b01111000100001111101101011111010;
		correct = 32'b10001011010101000111101110011000;
		#400 //-902.09155 * 2.2043795e+34 = -4.0922696e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110101011011110011010110001110;
		b = 32'b10101001100110000111100100011000;
		correct = 32'b11001011010010001101000001111100;
		#400 //8.911237e-07 * -6.7711624e-14 = -13160572.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001101100100010110000001000111;
		b = 32'b10100001010011011101001000010101;
		correct = 32'b00101011101101001101000110101001;
		#400 //-8.959493e-31 * -6.9734743e-19 = 1.2847962e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110011010111100100010111111001;
		b = 32'b11111111111110111000110100101000;
		correct = 32'b11111111111110111000110100101000;
		#400 //-5.1752043e-08 * nan = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001111011011111110110011010110;
		b = 32'b00111100100010110000101100010101;
		correct = 32'b10010010010111001101111010010110;
		#400 //-1.1829223e-29 * 0.016973058 = -6.969412e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101011111011100000001010010100;
		b = 32'b10100011000100011111111010110001;
		correct = 32'b01001000010100001010110001110110;
		#400 //-1.6911633e-12 * -7.914399e-18 = 213681.84
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000110010000011001001010000011;
		b = 32'b11100111111100010110001100001111;
		correct = 32'b10011101110011010100101001110000;
		#400 //12388.628 * -2.2798353e+24 = -5.4340015e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001000011001100010001011101111;
		b = 32'b10010101010000011101010010011101;
		correct = 32'b01110010100101111111100110110010;
		#400 //-235659.73 * -3.9143762e-26 = 6.020365e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100110011000001101101101011111;
		b = 32'b11001101010110000000101000111101;
		correct = 32'b10011000100001010011100101010000;
		#400 //7.8012915e-16 * -226534350.0 = -3.4437565e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111011101010011100000111101010;
		b = 32'b01111101110111010110010001001101;
		correct = 32'b10111101010001000100101101001101;
		#400 //-1.7628624e+36 * 3.6785022e+37 = -0.047923375
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010111111101000011100000010100;
		b = 32'b01010110111101101000101001000011;
		correct = 32'b01000000011111011001011100000100;
		#400 //537043380000000.0 * 135536845000000.0 = 3.9623423
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110101111101011100110001100011;
		b = 32'b11010110101110110011011011010111;
		correct = 32'b10011110101010000000110111110100;
		#400 //1.8313407e-06 * -102922105000000.0 = -1.7793463e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110001001000001110101100010011;
		b = 32'b11110100111111001011000100101111;
		correct = 32'b10111011101000110000011001010111;
		#400 //7.968286e+29 * -1.6016266e+32 = -0.004975121
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101110110011010111000100100100;
		b = 32'b01110100110101111011001000101010;
		correct = 32'b10111001011100111101010001111010;
		#400 //-3.1790603e+28 * 1.3671355e+32 = -0.0002325344
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110101000000010111111010011100;
		b = 32'b11010100011010011100100011011111;
		correct = 32'b01100000000011011100110010111110;
		#400 //-1.6415387e+32 * -4016389800000.0 = 4.0871002e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111000011001111011110011001;
		b = 32'b00001010100110001001100000001001;
		correct = 32'b11101011111011000111111010010000;
		#400 //-8.402299e-06 * 1.4694257e-32 = -5.7180834e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110011000000001001100100101;
		b = 32'b11001011010010101100000001110010;
		correct = 32'b10110010100011010111011000100111;
		#400 //0.21882303 * -13287538.0 = -1.646829e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101110110110110001001010111001;
		b = 32'b10111100100001101100010100110010;
		correct = 32'b00110001110100000001000101011101;
		#400 //-9.962293e-11 * -0.016451452 = 6.0555707e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100111110011111010111100000111;
		b = 32'b10101011010011001101111100100111;
		correct = 32'b10111100000000011100000111000100;
		#400 //5.7643807e-15 * -7.2785045e-13 = -0.0079197325
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001000010101111010101111010111;
		b = 32'b10010011000111100100111101101011;
		correct = 32'b10110100101011100110000011101110;
		#400 //6.4901206e-34 * -1.998156e-27 = -3.248055e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111000010110000010011001100100;
		b = 32'b11001010100101111001110100111001;
		correct = 32'b01101101001101100111101111111000;
		#400 //-1.7536168e+34 * -4968092.5 = 3.5297588e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010100001101111110101001110;
		b = 32'b01100011011101001100010010010101;
		correct = 32'b10010110100011010010111100011001;
		#400 //-0.0010298879 * 4.5151708e+21 = -2.2809501e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111111111100010110001100110101;
		b = 32'b00000111101110100100000000110101;
		correct = 32'b01111111111100010110001100110101;
		#400 //nan * 2.8023907e-34 = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011100011000101010001111010010;
		b = 32'b10100101000101001101101101100101;
		correct = 32'b00110110110000101110001001101001;
		#400 //-7.498886e-22 * -1.2911287e-16 = 5.808008e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101011011111111111010001100101;
		b = 32'b10111100011101110000110001111101;
		correct = 32'b00101110100001001001110101000010;
		#400 //-9.0933364e-13 * -0.015078661 = 6.0305996e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101011111010100101111011100101;
		b = 32'b01001100011000111111110100110000;
		correct = 32'b00011111000000111001010100110111;
		#400 //1.6653039e-12 * 59765950.0 = 2.7863757e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101011010011011110000010011101;
		b = 32'b00110000011010011111010010101001;
		correct = 32'b01111010011000010100011010101010;
		#400 //2.488905e+26 * 8.511259e-10 = 2.92425e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101011100110110001000011010110;
		b = 32'b11010010100100101101010010001010;
		correct = 32'b00011000100001110010110111101011;
		#400 //-1.1018085e-12 * -315315520000.0 = 3.4943047e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001110110101101110101101001010;
		b = 32'b00001111001110000101111101000010;
		correct = 32'b10111111000101010011010100001011;
		#400 //-5.298165e-30 * 9.0902464e-30 = -0.5828406
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010000000010110110111111101110;
		b = 32'b10010100011010011111100001000011;
		correct = 32'b11111011000110001001000100000001;
		#400 //9357474000.0 * -1.1812455e-26 = -7.9217015e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101001101110101001011101111001;
		b = 32'b11001001101111111110111100011100;
		correct = 32'b11011111011110001101111111011100;
		#400 //2.819694e+25 * -1572323.5 = -1.7933294e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010000001001101101001011010111;
		b = 32'b00010111100100110010111010111100;
		correct = 32'b01111000000100010001010011001001;
		#400 //11195342000.0 * 9.51145e-25 = 1.1770385e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101001000000101101111011000111;
		b = 32'b00101001111101011001110111000110;
		correct = 32'b10111110100010000110011100100101;
		#400 //-2.9059027e-14 * 1.0907555e-13 = -0.26641193
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100011000001110110101000110100;
		b = 32'b01101101011010101001000100100010;
		correct = 32'b10110101000100111100100111000010;
		#400 //-2.4979632e+21 * 4.5371842e+27 = -5.5055364e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001001011000111011001000010110;
		b = 32'b10001100101110100011111110111000;
		correct = 32'b00111100000111000111110000000000;
		#400 //-2.7407867e-33 * -2.8696187e-31 = 0.009551048
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011111000000001000111000110001;
		b = 32'b00100110101100000001110000100100;
		correct = 32'b00110111101110101101111101111101;
		#400 //2.7222672e-20 * 1.2220081e-15 = 2.2276998e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011111010111011101001111011111;
		b = 32'b10111110010001111011101100100111;
		correct = 32'b01100000100011100010100100101101;
		#400 //-1.5984365e+19 * -0.19504987 = 8.195015e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010011011111011100110000011110;
		b = 32'b10111011100001001011100011110010;
		correct = 32'b01010111011101001100010001010010;
		#400 //-1090051240000.0 * -0.0040503675 = 269124030000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011101101011001011011011101010;
		b = 32'b01101101101010100110010010001000;
		correct = 32'b00101111100000011011111010000001;
		#400 //1.555674e+18 * 6.5917483e+27 = 2.3600324e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010100000100110100000101001111;
		b = 32'b00111001000101111011111000001000;
		correct = 32'b11011010011110000110111000000110;
		#400 //-2529823600000.0 * 0.00014471274 = -1.7481692e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100000100001011001110111000111;
		b = 32'b10111010000000111111101110101001;
		correct = 32'b10100110000000011001010110000000;
		#400 //2.2635485e-19 * -0.00050347537 = -4.4958476e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100110000100110000110001111010;
		b = 32'b01010001011011101000000101101001;
		correct = 32'b00010100000111011101010110110111;
		#400 //5.101778e-16 * 64023335000.0 = 7.968622e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010000100111011001010011100001;
		b = 32'b00101011101011110010000011000010;
		correct = 32'b00100100011001100101100111010011;
		#400 //6.2154965e-29 * 1.244359e-12 = 4.9949384e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001110110001110110111000110010;
		b = 32'b10010010110011110101000111000100;
		correct = 32'b10111011011101100100001000110111;
		#400 //4.91634e-30 * -1.3083693e-27 = -0.0037576088
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011000000101110000001100001111;
		b = 32'b00001110011011000100100011000100;
		correct = 32'b11001001001000111001110011001110;
		#400 //-1.9517837e-24 * 2.9124281e-30 = -670156.9
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110101110110111011101100000000;
		b = 32'b01110010111000100000101010010110;
		correct = 32'b10000010011110001101101001001010;
		#400 //-1.6371196e-06 * 8.9544205e+30 = -1.8282808e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111100110000001111010111011010;
		b = 32'b01001101110100100010100011000111;
		correct = 32'b00101110011010110000110010110001;
		#400 //0.023554731 * 440735970.0 = 5.3444086e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101010001011000110111000001001;
		b = 32'b10110100110100001110000000111101;
		correct = 32'b00110100110100110101010011010100;
		#400 //-1.5314845e-13 * -3.8906174e-07 = 3.9363533e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111110001010100110110000111100;
		b = 32'b11101110001111110010001101001111;
		correct = 32'b11001111011001000100000101011000;
		#400 //5.6632686e+37 * -1.478858e+28 = -3829487600.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001111110101000001101101010000;
		b = 32'b11100011000101101111011110011011;
		correct = 32'b00101100001100111101011010001110;
		#400 //-7117119500.0 * -2.7848535e+21 = 2.5556532e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111101101101111001110111101;
		b = 32'b10100000001010001100100010001100;
		correct = 32'b11100111000010101011111010111111;
		#400 //93671.48 * -1.4296509e-19 = -6.552052e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011100010111111110010001010101;
		b = 32'b10001100010100110111110101000100;
		correct = 32'b01001111100001111000000110100110;
		#400 //-7.4079623e-22 * -1.6292544e-31 = 4546841600.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001000110001011101111101011010;
		b = 32'b01111011010001111011011100110001;
		correct = 32'b00001100111111011010001100101111;
		#400 //405242.8 * 1.0369826e+36 = 3.9079035e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000101001011000110111001010101;
		b = 32'b00100000110001001110011000110101;
		correct = 32'b10100011111000000010111111111010;
		#400 //-8.107666e-36 * 3.335603e-19 = -2.4306448e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110010011010111011100001000110;
		b = 32'b01010101111000110001000100110001;
		correct = 32'b00011100000001001110000010101010;
		#400 //1.3720699e-08 * 31207872000000.0 = 4.396551e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001100010100010010111001101111;
		b = 32'b01000111011101100110101011000100;
		correct = 32'b01000100010110010101000011110111;
		#400 //54835644.0 * 63082.766 = 869.2651
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110110111101011010000011011101;
		b = 32'b10101101110001101000111001010000;
		correct = 32'b11001000100111100101100001110010;
		#400 //7.320296e-06 * -2.2573193e-11 = -324291.56
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111011001100001010001000101110;
		b = 32'b00101010110110010000011110111110;
		correct = 32'b01001111110100000101100110000100;
		#400 //0.0026952135 * 3.8552316e-13 = 6991055000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110011001001011010001111111111;
		b = 32'b11101000001011001001101111100011;
		correct = 32'b11001010011101011010101001000110;
		#400 //1.3123401e+31 * -3.2604905e+24 = -4024977.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011011000010110100000101100100;
		b = 32'b01001111111010000000111011001001;
		correct = 32'b10001010100110011001111101111000;
		#400 //-1.1518939e-22 * 7786566000.0 = -1.479335e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000100011001100111011011101110;
		b = 32'b10100111010010100011010101100011;
		correct = 32'b00011100100100011110001011100111;
		#400 //-2.709098e-36 * -2.8062072e-15 = 9.653948e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001001011010111011111110011000;
		b = 32'b10000011111010000001110000011100;
		correct = 32'b11000101000000100000000110101110;
		#400 //2.8377183e-33 * -1.3642188e-36 = -2080.105
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100100100010101001000011011111;
		b = 32'b01011111000000001011001000101100;
		correct = 32'b10000101000010011101000100001001;
		#400 //-6.009338e-17 * 9.273523e+18 = -6.480103e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100001010101110001001101000001;
		b = 32'b00101111110100010010010101000111;
		correct = 32'b10110001000000111010000100000110;
		#400 //-7.2870316e-19 * 3.8043366e-10 = -1.915454e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110100101101000010000000011101;
		b = 32'b00111010000011011100010001000101;
		correct = 32'b11111010001000101010001001000010;
		#400 //-1.1416806e+32 * 0.00054079696 = -2.1111077e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011110100111010111110101000110;
		b = 32'b01010011000000110011001100010010;
		correct = 32'b11001011000110011010011000010100;
		#400 //-5.674152e+18 * 563497530000.0 = -10069524.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101111011000100111010111111111;
		b = 32'b01100011001010111000011111101100;
		correct = 32'b11001011101010001111110101101010;
		#400 //-7.008626e+28 * 3.1641874e+21 = -22149844.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011011010001101110011011110101;
		b = 32'b11001100001111110101011101010100;
		correct = 32'b11001110100001010000111011011101;
		#400 //5.5985985e+16 * -50158930.0 = -1116171900.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011101001001001011111111110;
		b = 32'b00111000110011111001000000001100;
		correct = 32'b11010010010010110000000011110010;
		#400 //-21573628.0 * 9.89736e-05 = -217973560000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000011000000001011011000111011;
		b = 32'b01010111000110000000011000110111;
		correct = 32'b10101011010110001011111001000011;
		#400 //-128.71184 * 167152460000000.0 = -7.7002657e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000011111000011000111011100111;
		b = 32'b10000110001011001110011111111100;
		correct = 32'b00111101001001101111101001000000;
		#400 //-1.325712e-36 * -3.252004e-35 = 0.040766
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110010000101110101001111001010;
		b = 32'b11111001111001001000110100011000;
		correct = 32'b00110111101010011000000001101010;
		#400 //-2.997346e+30 * -1.4833818e+35 = 2.0206167e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011100010011000100100110111110;
		b = 32'b11001000110111010010111110011011;
		correct = 32'b10010010111011000111000101000010;
		#400 //6.759325e-22 * -452988.84 = -1.4921614e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111110100001110000110010000101;
		b = 32'b11101100010111001011101011101010;
		correct = 32'b01010001100111001010000011000101;
		#400 //-8.975539e+37 * -1.0673854e+27 = 84089020000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000110101100000101010001001110;
		b = 32'b11010010001010011111000111100101;
		correct = 32'b10110100000001001100111100000100;
		#400 //22570.152 * -182476950000.0 = -1.236877e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010010100010010110011111010101;
		b = 32'b10010000110111011010010010101001;
		correct = 32'b11000001000111101011010001101011;
		#400 //8.671512e-28 * -8.742283e-29 = -9.919047
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111111011101000110011101010010;
		b = 32'b10010101010100011000001101110001;
		correct = 32'b11101001100101010101000011010110;
		#400 //0.95470154 * -4.2310903e-26 = -2.256396e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111011111000001011110110111010;
		b = 32'b01001101101001001101110101010100;
		correct = 32'b01101101101011100111110011100100;
		#400 //2.3338452e+36 * 345746050.0 = 6.750172e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110001011111010101000010111011;
		b = 32'b00110011010011010011101101001111;
		correct = 32'b01111101100111011111110100110101;
		#400 //1.2543569e+30 * 4.7784223e-08 = 2.625044e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001001001010101000000010010001;
		b = 32'b01110001101010000010011111110010;
		correct = 32'b10010111000000011100100100110001;
		#400 //-698377.06 * 1.6653367e+30 = -4.1936087e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011110000110011000011011101111;
		b = 32'b01110010110101001101010011010001;
		correct = 32'b10101010101110001010101011000101;
		#400 //-2.765698e+18 * 8.431117e+30 = -3.280346e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000110001011001110010010000100;
		b = 32'b00001101100100101010001100011001;
		correct = 32'b11111000000101101110101100100110;
		#400 //-11065.129 * 9.037209e-31 = -1.2243967e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101101100001101110100001010100;
		b = 32'b11000100011100101101001000100111;
		correct = 32'b01101000100011100011101011001001;
		#400 //-5.2189823e+27 * -971.2836 = 5.3732835e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010101010011100111101110000111;
		b = 32'b11001000011010010111110000011011;
		correct = 32'b00001100011000100110010011010101;
		#400 //-4.1698815e-26 * -239088.42 = 1.744075e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101000010001110010010100010010;
		b = 32'b10100110110101110111100011111010;
		correct = 32'b01000000111011001001100111101001;
		#400 //-1.10547574e-14 * -1.4951413e-15 = 7.393788
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101010110100010001011101001010;
		b = 32'b11101010011001001100010101100101;
		correct = 32'b10111111111010011111101000111111;
		#400 //1.2638774e+26 * -6.9141814e+25 = -1.8279494
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010101010110110010101101101111;
		b = 32'b11000100111011101011101000111000;
		correct = 32'b11001111111010110000011011110110;
		#400 //15061225000000.0 * -1909.8193 = -7886204000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100101011101111100001110000100;
		b = 32'b10101101011010101000101100111010;
		correct = 32'b11110111100001110011011011110001;
		#400 //7.3126947e+22 * -1.33322745e-11 = -5.4849564e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010101100001101001001001101111;
		b = 32'b00111011110000101011010000010011;
		correct = 32'b01011001001100001111000000100001;
		#400 //18495436000000.0 * 0.0059418767 = 3112726300000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000101110010000001000000011010;
		b = 32'b11101100010011111111101011111001;
		correct = 32'b10011000111101100100000100100111;
		#400 //6402.0127 * -1.0057313e+27 = -6.3655297e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111011101111011001000110101001;
		b = 32'b01011001111110001000001001010001;
		correct = 32'b10100001010000110100100010000101;
		#400 //-0.0057851863 * 8743635000000000.0 = -6.616455e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001001110100110010111001100000;
		b = 32'b01110011100001110011011111101111;
		correct = 32'b00010101110001111110100001010001;
		#400 //1729996.0 * 2.1426225e+31 = 8.074199e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001100000000011011101101101011;
		b = 32'b00110000001001001101101011001100;
		correct = 32'b00011011010010010111010101110001;
		#400 //9.994198e-32 * 5.997378e-10 = 1.6664278e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101011110011000001111001000100;
		b = 32'b10000100001111110110110011110111;
		correct = 32'b11100111000010000111110010110011;
		#400 //1.4503472e-12 * -2.2501976e-36 = -6.4454214e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011010111010011011001110011100;
		b = 32'b00100111010100010011101101110110;
		correct = 32'b11110011000011101111100000101000;
		#400 //-3.2890576e+16 * 2.903681e-15 = -1.13272e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101111011100100100100000011000;
		b = 32'b01001110101011011001001000001100;
		correct = 32'b11100000001100101010101111010011;
		#400 //-7.498253e+28 * 1456014800.0 = -5.1498464e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000101101001110100110110110000;
		b = 32'b00100111011100010100010010100110;
		correct = 32'b10011101101100011000010011011111;
		#400 //-1.5733142e-35 * 3.3482683e-15 = -4.6988895e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011010111110110000010001011001;
		b = 32'b01101101010000110001001101001001;
		correct = 32'b00101101001001001011010011011101;
		#400 //3.53275e+16 * 3.7733057e+27 = 9.36248e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010110001101111110110011011101;
		b = 32'b00110111111101111001000011011010;
		correct = 32'b11011101101111100011000011111000;
		#400 //-50556987000000.0 * 2.9512146e-05 = -1.7130908e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101001111111100010010110100100;
		b = 32'b00110001001010100010011101111111;
		correct = 32'b01111000001111110010111100101100;
		#400 //3.8405614e+25 * 2.4760707e-09 = 1.551071e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110011101101100101001001010011;
		b = 32'b11011010101100101000011001101001;
		correct = 32'b10011000100000101011100011011001;
		#400 //8.49001e-08 * -2.5125166e+16 = -3.379086e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110011101110010010011010110001;
		b = 32'b01000101010101100010100010011000;
		correct = 32'b10101101110111010101001101000001;
		#400 //-8.621772e-08 * 3426.537 = -2.5161763e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110101010000010000000011001110;
		b = 32'b01101111011010000101110010100100;
		correct = 32'b11000101010101001010001100100111;
		#400 //-2.4466055e+32 * 7.191252e+28 = -3402.197
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101110100000110001010000001101;
		b = 32'b10011010001100111000101100000101;
		correct = 32'b01010011101110101110010110100000;
		#400 //-5.960752e-11 * -3.712863e-23 = 1605432800000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101100111111101100001010000000;
		b = 32'b11000011001010011011110100110011;
		correct = 32'b11101001010000000001110100101111;
		#400 //2.4638853e+27 * -169.73906 = -1.4515723e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001100111111000100000001011111;
		b = 32'b11000111101101100101110100101110;
		correct = 32'b11000100101100010000110110110100;
		#400 //132252410.0 * -93370.36 = -1416.4282
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000001111101101111010000001101;
		b = 32'b10100000010001100000100001010010;
		correct = 32'b11100001000111111001111011010010;
		#400 //30.869165 * -1.6774005e-19 = -1.8402978e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010000110111111110001111110111;
		b = 32'b10101001101000011100100010101011;
		correct = 32'b11100110101100010010001100110001;
		#400 //30050073000.0 * -7.1846466e-14 = -4.18254e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011100110000100101000010001010;
		b = 32'b00101101111101111111011100010000;
		correct = 32'b01101110010010001001110001101110;
		#400 //4.375576e+17 * 2.8190367e-11 = 1.5521528e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000100100001110000000001001101;
		b = 32'b11110011001111011011011100101110;
		correct = 32'b00010000101101100010101101000111;
		#400 //-1080.0094 * -1.5030814e+31 = 7.185302e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110110100010011110101101101010;
		b = 32'b11011001110011000100011111110010;
		correct = 32'b11011100001011001101011001100011;
		#400 //1.3986708e+33 * -7187500000000000.0 = -1.9459767e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100011000000001100010010101000;
		b = 32'b11001011000001011011111100000000;
		correct = 32'b00010111011101100111100011010000;
		#400 //-6.9805375e-18 * -8765184.0 = 7.9639374e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100011011111001100001101000100;
		b = 32'b11001101011101101110111101010100;
		correct = 32'b10010101100000110000010101011011;
		#400 //1.37022965e-17 * -258929980.0 = -5.291893e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011001110010100011110100110101;
		b = 32'b11100010010110011110111101101000;
		correct = 32'b00110110111011011000111111111010;
		#400 //-7115655400000000.0 * -1.0050486e+21 = 7.0799115e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110001101110011100011000101000;
		b = 32'b00110011001000111001100101010101;
		correct = 32'b10111110000100010101100110001110;
		#400 //-5.4067364e-09 * 3.809085e-08 = -0.14194319
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110001100010000100111111000000;
		b = 32'b00111100110010101111010011011011;
		correct = 32'b11110100001010111110111111100111;
		#400 //-1.349964e+30 * 0.02477496 = -5.448905e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111001011011101110101111101010;
		b = 32'b11001101000111101000100000011000;
		correct = 32'b01101011110000001110100001011010;
		#400 //-7.753447e+34 * -166232450.0 = 4.66422e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100010010000111101010000100010;
		b = 32'b01010001110000111110110000000101;
		correct = 32'b01001111111111111110000011001010;
		#400 //9.031002e+20 * 105184800000.0 = 8585843700.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110101111100110111101010001001;
		b = 32'b01000111010011010000011001001100;
		correct = 32'b01101110000110000000000111101001;
		#400 //6.1729172e+32 * 52486.297 = 1.1761008e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111111011010010000101101000;
		b = 32'b01001010011111100011111010111000;
		correct = 32'b10101100111011101100010001110010;
		#400 //-2.8268158e-05 * 4165550.0 = -6.7861767e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010110010110110101101100010110;
		b = 32'b00000001100000101010111000111100;
		correct = 32'b11010100010101101101101100110011;
		#400 //-1.7719421e-25 * 4.800447e-38 = -3691202200000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100001001111010111011100010010;
		b = 32'b00111111000011100110100000111110;
		correct = 32'b11100001101010100100110000010000;
		#400 //-2.1843841e+20 * 0.5562781 = -3.9267842e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011101001010111111000011010011;
		b = 32'b01011001011001101111110010100000;
		correct = 32'b00000011001111101000111101010101;
		#400 //2.2756165e-21 * 4063563000000000.0 = 5.600052e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011111010010100101010100010101;
		b = 32'b00010100011111110110111011010010;
		correct = 32'b11001010010010101100100000010101;
		#400 //-4.2845542e-20 * 1.28960654e-26 = -3322373.2
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100011011101100110000100101011;
		b = 32'b01001001111110100011111000111111;
		correct = 32'b00011000111111000000110000101011;
		#400 //1.3356263e-17 * 2049991.9 = 6.515276e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100001110010110101010110011100;
		b = 32'b10101101011000110010101101000011;
		correct = 32'b10110011111001010010001111110110;
		#400 //1.3778476e-18 * -1.2913062e-11 = -1.0670185e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011000111001100100111100101101;
		b = 32'b00110001111011001101010101000000;
		correct = 32'b00100110011110001111001011000100;
		#400 //5.9533554e-24 * 6.8927477e-09 = 8.6371293e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100011101100011101000101001000;
		b = 32'b10010000010000011011100101011000;
		correct = 32'b01010010111010101111101011100111;
		#400 //-1.9279013e-17 * -3.8205322e-29 = 504615900000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100110101001000100011011111000;
		b = 32'b10111111110011111100100110010101;
		correct = 32'b01100110010010100110010011101010;
		#400 //-3.8788862e+23 * -1.6233393 = 2.389449e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010001011111101110001111111111;
		b = 32'b00001001110001111001100110101110;
		correct = 32'b01000111001000110111010011100111;
		#400 //2.0107324e-28 * 4.8052027e-33 = 41844.902
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111110111100010100100100001011;
		b = 32'b01011111110111001110011101001011;
		correct = 32'b10011110100010111100111101011110;
		#400 //-0.4712604 * 3.1835548e+19 = -1.4802963e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010010110100110100100111100111;
		b = 32'b11101110001100100100000110111100;
		correct = 32'b10100100000101111011100000010101;
		#400 //453739000000.0 * -1.379195e+28 = -3.289883e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001001111010101101010101010001;
		b = 32'b11001011111011110101001100011101;
		correct = 32'b10111101011110110011001000010111;
		#400 //1923754.1 * -31368762.0 = -0.061327066
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100111100000100011011000111011;
		b = 32'b11111000010000001001110110000011;
		correct = 32'b00101110101011010000111110101010;
		#400 //-1.229816e+24 * -1.5626808e+34 = 7.869912e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001101001011101111010010111000;
		b = 32'b00010101010011101111010111011110;
		correct = 32'b10110111010110000110100101111001;
		#400 //-5.391246e-31 * 4.1795324e-26 = -1.28991605e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111111101111101001001110101111;
		b = 32'b10000111100100101101010111001110;
		correct = 32'b11110111101001100010000101111011;
		#400 //1.488882 * -2.2093302e-34 = -6.739065e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110001011001101010111010111110;
		b = 32'b01010110111110010110110111000000;
		correct = 32'b01011001111011001100001010010000;
		#400 //1.14228484e+30 * 137124880000000.0 = 8330252300000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001110000101011001110000101111;
		b = 32'b10110101111101011010110000011010;
		correct = 32'b01010111100110111110011001000101;
		#400 //-627510200.0 * -1.8304011e-06 = 342826600000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010110111100000111000101011100;
		b = 32'b11000110011100100010010111011000;
		correct = 32'b10001111111111100011001010001100;
		#400 //3.884563e-25 * -15497.461 = -2.5065804e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100011111000001110101000101111;
		b = 32'b01111001100010010100100111000100;
		correct = 32'b10101001110100011011001011000100;
		#400 //-8.297891e+21 * 8.91051e+34 = -9.3124754e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000001110110000011001011101001;
		b = 32'b01100101111101110000111000011110;
		correct = 32'b10011011011000000000011011001100;
		#400 //-27.024858 * 1.4583562e+23 = -1.8531042e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010000101000001011111100011111;
		b = 32'b01001110001010100101011010001011;
		correct = 32'b00000001111100011001010111000011;
		#400 //6.340334e-29 * 714449600.0 = 8.8744316e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111111110001101110100000001010;
		b = 32'b00110010001011001111101100000001;
		correct = 32'b01111111110001101110100000001010;
		#400 //nan * 1.0068789e-08 = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110110011000011001011100100;
		b = 32'b01011000001000101101101100101000;
		correct = 32'b10011110001000000111111010000000;
		#400 //-6.085598e-06 * 716248600000000.0 = -8.496489e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111000101100001100110010110111;
		b = 32'b01011000000010001110001000100100;
		correct = 32'b01100000001001010101001101101011;
		#400 //2.8687386e+34 * 602019400000000.0 = 4.7651932e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111001111111110011110111111100;
		b = 32'b00100110100100100011101001011010;
		correct = 32'b11010010110111110110110011010100;
		#400 //-0.00048683572 * 1.0146601e-15 = -479801770000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110100100000000100110011000011;
		b = 32'b11000111010100100101001101110011;
		correct = 32'b11101100100111000010100101000110;
		#400 //8.131969e+31 * -53843.45 = -1.5102987e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010001000110111011001010000011;
		b = 32'b00110000011101110011110000100010;
		correct = 32'b00100000001000010011011110011001;
		#400 //1.2282352e-28 * 8.994353e-10 = 1.3655626e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011000010010111100101011001110;
		b = 32'b00010011010011000100001101111101;
		correct = 32'b01000100011111110110100011000000;
		#400 //2.6339525e-24 * 2.5781694e-27 = 1021.6367
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000011110010000100001110110001;
		b = 32'b10110001110010110001110110001101;
		correct = 32'b11010001011111000110100000011100;
		#400 //400.52884 * -5.911437e-09 = -67754900000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100010001100000101110011100111;
		b = 32'b00010011011111010010010001100110;
		correct = 32'b11001110001100100101101010011011;
		#400 //-2.390163e-18 * 3.1951035e-27 = -748070600.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001110100011000011100011011100;
		b = 32'b11011100011001101110011101111010;
		correct = 32'b10110001100110110111011001001110;
		#400 //1176268300.0 * -2.5997502e+17 = -4.5245434e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111010000101110000000110101111;
		b = 32'b10001001000010001000001010110010;
		correct = 32'b11110000100011011001011110100010;
		#400 //0.0005760444 * -1.6431857e-33 = -3.505656e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001000011111110010100101101000;
		b = 32'b10101111110101011111110001101011;
		correct = 32'b10011000000110001010000101001101;
		#400 //7.6784944e-34 * -3.8923828e-10 = -1.9726976e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001000101100001010001111001110;
		b = 32'b11001111000001111110111111011100;
		correct = 32'b10111001001001100101001110001110;
		#400 //361758.44 * -2280643600.0 = -0.0001586212
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011000001011111111000010110011;
		b = 32'b00000000111101100011100100000100;
		correct = 32'b01010110101101101110110100111010;
		#400 //2.2739742e-24 * 2.2611985e-38 = 100565000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100111011100111011111101111100;
		b = 32'b10101011101100101101001111010100;
		correct = 32'b00111011001011100111011111101010;
		#400 //-3.3826828e-15 * -1.2706455e-12 = 0.0026621767
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001001000000100001111011111110;
		b = 32'b11101100000001010000010111010101;
		correct = 32'b10011100011110100110101001101011;
		#400 //532975.9 * -6.432587e+26 = -8.2855603e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001101101001010110110100101000;
		b = 32'b00100110001110001000000111110110;
		correct = 32'b11100110111001011000011001110011;
		#400 //-346924300.0 * 6.4013954e-16 = -5.4195104e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011010110101001111100011111101;
		b = 32'b00110101100101110010101111011000;
		correct = 32'b00100100101101000101010000011011;
		#400 //8.808341e-23 * 1.1263137e-06 = 7.8205037e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110100100101001110111011000010;
		b = 32'b00011001001110011110101101100000;
		correct = 32'b01011010110011010001001001000111;
		#400 //2.7740867e-07 * 9.6118094e-24 = 2.8861233e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001011101001011010001111000000;
		b = 32'b01100000011011100010101000000001;
		correct = 32'b00101010101100100000101101010101;
		#400 //21710720.0 * 6.864612e+19 = 3.1627015e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001001000100010001001001101011;
		b = 32'b01100011111101000110010001110011;
		correct = 32'b00100100100101111111011001010111;
		#400 //594214.7 * 9.0164874e+21 = 6.590313e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111111000111001010101101000101;
		b = 32'b11110010000110111101110000101101;
		correct = 32'b10001100100000001010101000010011;
		#400 //0.61198837 * -3.0871266e+30 = -1.9823882e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111011011111111010011000110000;
		b = 32'b11100010100000011110010101110010;
		correct = 32'b01011000011110111110101011001000;
		#400 //-1.3274064e+36 * -1.1980816e+21 = 1107943200000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011001001110010101010000110011;
		b = 32'b10000111000100100110111001110000;
		correct = 32'b01010001101000100000000001011111;
		#400 //-9.58128e-24 * -1.1016274e-34 = 86973870000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100101101110110010100101011111;
		b = 32'b01001110001000000111011100111100;
		correct = 32'b00010111000101010100101101110001;
		#400 //3.2467363e-16 * 673042200.0 = 4.8239717e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101001011010010101111110010100;
		b = 32'b01011011111010111101011100100100;
		correct = 32'b10001100111111010101001001110100;
		#400 //-5.1819294e-14 * 1.3276634e+17 = -3.9030447e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100000010111100010011101010011;
		b = 32'b10111100110000101010000000001011;
		correct = 32'b10100011000100100001101011010001;
		#400 //1.8817143e-19 * -0.023757955 = -7.9203545e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111011000011010001110111101001;
		b = 32'b10111011100001000001100001111110;
		correct = 32'b10111111000010001011110111010000;
		#400 //0.002153272 * -0.00403124 = -0.5341463
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010110010111001000110010110110;
		b = 32'b01011111111101101100011010001111;
		correct = 32'b10110101111001001100101100110001;
		#400 //-60624227000000.0 * 3.5564115e+19 = -1.704646e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100010110000000100001010101100;
		b = 32'b00101100111100110011010001011011;
		correct = 32'b00110101010010100110000000101011;
		#400 //5.2112296e-18 * 6.912288e-12 = 7.5390807e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110101110100011110010100101011;
		b = 32'b10101000011101001100110110100010;
		correct = 32'b11001100110110110111111011001101;
		#400 //1.563841e-06 * -1.358931e-14 = -115078760.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101011111001010110000101101011;
		b = 32'b01010001111011111100001001100000;
		correct = 32'b10011001011101001110101100010001;
		#400 //-1.6298468e-12 * 128719780000.0 = -1.2661976e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011100110101010110111101110011;
		b = 32'b11011000101101111101101100010110;
		correct = 32'b00000011100101001001011111011101;
		#400 //-1.4123967e-21 * -1617212800000000.0 = 8.733524e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010101101100011111010011101110;
		b = 32'b10101001010011100100010000110011;
		correct = 32'b10101011110111001101110101010001;
		#400 //7.187616e-26 * -4.5800342e-14 = -1.5693368e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110000010101101110011100100111;
		b = 32'b01101010000001101001111001011010;
		correct = 32'b01000101110011000101011001010001;
		#400 //2.6603695e+29 * 4.0685963e+25 = 6538.7896
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101011110000111111011001100110;
		b = 32'b01110011011010101011101110101100;
		correct = 32'b10110111110101011011011101111110;
		#400 //-4.7380824e+26 * 1.8597472e+31 = -2.5477024e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101010000010100110000110000001;
		b = 32'b00101010100100011000101010010110;
		correct = 32'b00111110111100110110011110110011;
		#400 //1.229069e-13 * 2.5853337e-13 = 0.47540054
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001111001000001011110011100000;
		b = 32'b00010111011100000110100001101000;
		correct = 32'b01110111001010110010100110101100;
		#400 //2696732700.0 * 7.767996e-25 = 3.4715936e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101010001010111011101100100111;
		b = 32'b11010101110011001110100101000100;
		correct = 32'b10010011110101101000110000011111;
		#400 //1.5252782e-13 * -28162780000000.0 = -5.4159365e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001010111001011000001000110000;
		b = 32'b00110110001101010001110101100111;
		correct = 32'b00010100001000100011001110010011;
		#400 //2.2100869e-32 * 2.6988216e-06 = 8.189081e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011000011010001000101010111011;
		b = 32'b01101101101100011111000110011010;
		correct = 32'b10101010001001110100011000100101;
		#400 //-1022730160000000.0 * 6.8838656e+27 = -1.4856916e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000000110110011010011010111111;
		b = 32'b10101111011100101000010110101000;
		correct = 32'b10010000111001011011111101000001;
		#400 //1.998812e-38 * -2.2057256e-10 = -9.0619247e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011110111000100000000111110010;
		b = 32'b01010011010011110110000000010101;
		correct = 32'b00001011000010111000000000100100;
		#400 //2.3929485e-20 * 890670200000.0 = 2.6866829e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000110110011010001100111100001;
		b = 32'b11110010000101100010001001110111;
		correct = 32'b10010100001011101101110011010111;
		#400 //26252.94 * -2.9737227e+30 = -8.828308e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001000011110010110010100110011;
		b = 32'b10101011111110111111011100001111;
		correct = 32'b11011011111111010110001110011011;
		#400 //255380.8 * -1.7903195e-12 = -1.4264537e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011010011000100101101111110110;
		b = 32'b10110100001100010101010010001110;
		correct = 32'b01100101101000110110001111010001;
		#400 //-1.5928614e+16 * -1.651517e-07 = 9.644838e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001110001100111111100010100100;
		b = 32'b11001010000111011101111101100010;
		correct = 32'b00000011100100011110101011001011;
		#400 //-2.218317e-30 * -2586584.5 = 8.57624e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010011111100011001110010010001;
		b = 32'b01000111110101101011000100000101;
		correct = 32'b00001011100100000000110011000101;
		#400 //6.099134e-27 * 109922.04 = 5.5485996e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000110000101000010011011001001;
		b = 32'b11001000011100000010001010110100;
		correct = 32'b00111101000111011111000001100110;
		#400 //-9481.696 * -245898.81 = 0.03855934
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010100111011011111101111110100;
		b = 32'b10111010110110100101110111111001;
		correct = 32'b00011001100010110111111110111011;
		#400 //-2.4030262e-26 * -0.0016660086 = 1.4423853e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010010101011101010010000110110;
		b = 32'b10011101001010000101001011111111;
		correct = 32'b11110101000001001100110111001010;
		#400 //375039660000.0 * -2.2277523e-21 = -1.683489e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010100001110101011110001111001;
		b = 32'b00111000010101011101111101001001;
		correct = 32'b11011011010111111000010011010100;
		#400 //-3208103900000.0 * 5.0991108e-05 = -6.2914966e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111101111010000011110110001001;
		b = 32'b01011101011100011001001010010111;
		correct = 32'b11011111111101100001110001000100;
		#400 //-3.858755e+37 * 1.08794635e+18 = -3.5468248e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011000000111110101100011011100;
		b = 32'b11010011111011101101101001011011;
		correct = 32'b00000011101010101100100101011000;
		#400 //-2.059513e-24 * -2051731200000.0 = 1.0037928e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010010011110001111001010101111;
		b = 32'b11001111011100110011111110110111;
		correct = 32'b01000010100000101111111110111001;
		#400 //-267305860000.0 * -4081039000.0 = 65.49946
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010111111101010000011001101011;
		b = 32'b00001001110101001100001101010001;
		correct = 32'b11001101100100110110100010111111;
		#400 //-1.5834374e-24 * 5.122082e-33 = -309139420.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001011011101101011001001101111;
		b = 32'b00001101000000111100010110011101;
		correct = 32'b00111101111011111010001010101001;
		#400 //4.7512115e-32 * 4.060536e-31 = 0.11700947
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100101101100011101101010101001;
		b = 32'b01100000011101011111010101100100;
		correct = 32'b11000100101110010001110101111100;
		#400 //-1.0498655e+23 * 7.0892727e+19 = -1480.9214
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110110101001010011010101111000;
		b = 32'b10011110100111000111000100100101;
		correct = 32'b11010111100001110010110001001011;
		#400 //4.923608e-06 * -1.6563938e-20 = -297248600000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000101010101101011000001111111;
		b = 32'b00110110010000010001100111000100;
		correct = 32'b00001110100011100100111101111100;
		#400 //1.0094649e-35 * 2.8774239e-06 = 3.5082243e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110101101011111001110100011111;
		b = 32'b01101100011110010001110111011000;
		correct = 32'b10001000101101000111011101011001;
		#400 //-1.3084244e-06 * 1.20465385e+27 = -1.0861414e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101001011100010000001101011011;
		b = 32'b01100011101011000010111110000111;
		correct = 32'b01000101001100110010101001001011;
		#400 //1.8210436e+25 * 6.3525294e+21 = 2866.6433
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110100111100101000110001010000;
		b = 32'b10110101011011100000100010100010;
		correct = 32'b10111111000000100110110101110100;
		#400 //4.5178103e-07 * -8.867447e-07 = -0.5094826
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011111011100001001001011101100;
		b = 32'b10101001010110000111110111111000;
		correct = 32'b00110101100011100011110100000000;
		#400 //-5.0943508e-20 * -4.8070895e-14 = 1.0597578e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000101101001100110000000111000;
		b = 32'b10111011110000001011111100110001;
		correct = 32'b01001001010111001111100110010101;
		#400 //-5324.0273 * -0.005882167 = 905113.3
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001110011101001110100011110001;
		b = 32'b11111000110100011101001001000110;
		correct = 32'b10010101000101010110011111010000;
		#400 //1027226700.0 * -3.4045465e+34 = -3.0172204e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100010011101011100001010110111;
		b = 32'b11100110100110111000111110100101;
		correct = 32'b10111011010010100011011111111001;
		#400 //1.13337075e+21 * -3.673083e+23 = -0.0030856116
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011101001000010011010110011110;
		b = 32'b10101101011110101000001001101101;
		correct = 32'b01101111001001001011111000100100;
		#400 //-7.260228e+17 * -1.4239815e-11 = 5.0985408e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001001110001101111010111011110;
		b = 32'b10011110001011110111001111010000;
		correct = 32'b11101011000100010010011001101101;
		#400 //1629883.8 * -9.288372e-21 = -1.754757e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101100110010100010101011100001;
		b = 32'b11010000010111100001100001111010;
		correct = 32'b00011011111010010000011110011100;
		#400 //-5.745946e-12 * -14904584000.0 = 3.8551534e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100101000100110111000100000101;
		b = 32'b01010111011000010001110001000000;
		correct = 32'b00001101001001111010110001100100;
		#400 //1.278851e-16 * 247511450000000.0 = 5.1668356e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101010101111010010000100100010;
		b = 32'b01001000001110001011001010110011;
		correct = 32'b01100010000000110001001000110000;
		#400 //1.1432172e+26 * 189130.8 = 6.044585e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011010011110000001110110010101;
		b = 32'b01100100101000000100001010011001;
		correct = 32'b10110101010001100010101110010101;
		#400 //-1.745958e+16 * 2.3650223e+22 = -7.382417e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110001100100011011110001111101;
		b = 32'b00110111111000000000001001100011;
		correct = 32'b11111001001001101000110001111111;
		#400 //-1.4433022e+30 * 2.6703992e-05 = -5.404818e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110010010001111110001111001100;
		b = 32'b01111100101111100001000000000111;
		correct = 32'b10110101000001101001111001000111;
		#400 //-3.959226e+30 * 7.894892e+36 = -5.0149214e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111111110000010001000101000100;
		b = 32'b01000101011111001101001100000010;
		correct = 32'b10111001110000110111111000011010;
		#400 //-1.5083394 * 4045.188 = -0.0003728725
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011111111111110100111110100100;
		b = 32'b00011110011111000100001010100010;
		correct = 32'b01000001000000011000110001001011;
		#400 //1.08128455e-19 * 1.3354548e-20 = 8.096751
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010110110101011000101001101011;
		b = 32'b01001110001100111011101011010001;
		correct = 32'b00001000000110000001010001011001;
		#400 //3.449936e-25 * 753841200.0 = 4.5764755e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110010011000000101110100001100;
		b = 32'b11001011010010111000100001100010;
		correct = 32'b01100110100011010001100110101011;
		#400 //-4.4439763e+30 * -13338722.0 = 3.331636e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101110100011011000100011101010;
		b = 32'b00111110110101011000110010001011;
		correct = 32'b01101111001010011010101110010110;
		#400 //2.1901453e+28 * 0.41708788 = 5.25104e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110011010100010101000000000100;
		b = 32'b11001101111010010101100011100010;
		correct = 32'b11100100111001011010000111010100;
		#400 //1.658345e+31 * -489364540.0 = -3.3887723e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011111100101110010110010101001;
		b = 32'b11110000001101101100001010100100;
		correct = 32'b00101110110100111100000110100001;
		#400 //-2.1786535e+19 * -2.2624631e+29 = 9.6295645e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100110010111010010111011000010;
		b = 32'b01111100000011110110000001101111;
		correct = 32'b00101001110001010111011000100110;
		#400 //2.6112638e+23 * 2.9778174e+36 = 8.769053e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110111010111101001010110010010;
		b = 32'b11111100111011110001000110110101;
		correct = 32'b10111001111011100101100011111110;
		#400 //4.514545e+33 * -9.930545e+36 = -0.00045461202
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000001011101101001001101101101;
		b = 32'b00101011011001101000000100100101;
		correct = 32'b01010101100010001110110010101101;
		#400 //15.410993 * 8.189164e-13 = 18818762000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010100001010000100011010110101;
		b = 32'b11010010111011001001100111011101;
		correct = 32'b01000000101101100001001010111101;
		#400 //-2890963000000.0 * -508096840000.0 = 5.6897874
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101101101000000110100001111110;
		b = 32'b10011001000101000001110000000001;
		correct = 32'b01010100000010101010000100000001;
		#400 //-1.8236298e-11 * -7.657076e-24 = 2381626700000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000010001000100110100001101110;
		b = 32'b10011101010010011001101100010101;
		correct = 32'b10100100010011100011100111110011;
		#400 //1.193185e-37 * -2.6682304e-21 = -4.4718214e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011101010100011101110100101101;
		b = 32'b01011000001000110011001010111000;
		correct = 32'b10000100101001001001100111100001;
		#400 //-2.7775265e-21 * 717752900000000.0 = -3.869753e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101100101000000111010000110101;
		b = 32'b11010110110101010100001101111000;
		correct = 32'b11010101010000001001101110010100;
		#400 //1.5518152e+27 * -117242880000000.0 = -13235902000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000110000101001111010100101011;
		b = 32'b11000011001010001100011111000011;
		correct = 32'b00000010011000011110111100001001;
		#400 //-2.8015827e-35 * -168.78032 = 1.6598989e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011110000110011111101111100010;
		b = 32'b10011101100110101110000001001110;
		correct = 32'b10111111111111101000011001101111;
		#400 //8.151841e-21 * -4.0995386e-21 = -1.9884776
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010001110101111010101110011010;
		b = 32'b00011101001101011000101111100000;
		correct = 32'b01110100000110000000111100101001;
		#400 //115787120000.0 * 2.4027464e-21 = 4.818949e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110001011010101100000100110;
		b = 32'b01001010011110101110011111101101;
		correct = 32'b00110011001100001101110100011001;
		#400 //0.16928157 * 4110843.2 = 4.117928e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001010000101011110001101010010;
		b = 32'b01011001100111011010100010000001;
		correct = 32'b00101111111100110110001000001000;
		#400 //2455764.5 * 5547105400000000.0 = 4.4271098e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001000111001011101111100110111;
		b = 32'b01111001110001001111001011111001;
		correct = 32'b00001110100101010110010110100010;
		#400 //470777.72 * 1.2782728e+35 = 3.6829205e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100010100101101000010010110010;
		b = 32'b10011110111011111101001100101010;
		correct = 32'b11000011001000001010101110001111;
		#400 //4.079808e-18 * -2.5392445e-20 = -160.67015
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101011111110110010101001001000;
		b = 32'b11100101101000001110010001010101;
		correct = 32'b01000101110001111101000101111000;
		#400 //-6.072801e+26 * -9.497383e+22 = 6394.1836
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110001101011001110001110000110;
		b = 32'b10110101110100010111000101101101;
		correct = 32'b10111011010100110101000111110000;
		#400 //5.0317253e-09 * -1.5604725e-06 = -0.0032244883
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111100000001001010110101110110;
		b = 32'b01001001111000111111011101010010;
		correct = 32'b11110001100101001111111001010100;
		#400 //-2.7556056e+36 * 1867498.2 = -1.4755598e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000000111001111111110101111100;
		b = 32'b10110100100110010010111001011100;
		correct = 32'b00001011110000011101101010010101;
		#400 //-2.1304933e-38 * -2.8532202e-07 = 7.466978e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010010000100011110001001001001;
		b = 32'b01011010011100111000100111010011;
		correct = 32'b00110111000110010101100101000010;
		#400 //156641670000.0 * 1.713749e+16 = 9.140293e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100000000111101111001011001101;
		b = 32'b00110111001100010000001110000001;
		correct = 32'b10101000011001011101111110101110;
		#400 //-1.3463457e-19 * 1.0550838e-05 = -1.27605564e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010011110010101000011101111000;
		b = 32'b11100111001111110010111000100100;
		correct = 32'b10101100000001111001100100110001;
		#400 //1739712400000.0 * -9.0282314e+23 = -1.9269692e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100000000100101011001101111110;
		b = 32'b11000101001110111001011001011110;
		correct = 32'b11011010010010000011001111100010;
		#400 //4.2283725e+19 * -3001.398 = -1.408801e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010111100111110110101001000100;
		b = 32'b00110111100110111011100000101001;
		correct = 32'b00011111100000110000100110110001;
		#400 //1.0301959e-24 * 1.8563196e-05 = 5.549669e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001010010111001101100000101110;
		b = 32'b00101110110100011000110001011001;
		correct = 32'b10011011000001101110011001110001;
		#400 //-1.06332736e-32 * 9.5291504e-11 = -1.115868e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110000001001010110101101011;
		b = 32'b11001111100100110110000101011111;
		correct = 32'b00100101111001100111011000000001;
		#400 //-1.9770475e-06 * -4945264000.0 = 3.9978603e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101101000010000001000101111111;
		b = 32'b01110000111001000111000011100110;
		correct = 32'b00111011100110000111101111001010;
		#400 //2.6319446e+27 * 5.6559254e+29 = 0.0046534287
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001101000100010010001010000100;
		b = 32'b01111101001100000110001111011011;
		correct = 32'b00001111010100101010001101101101;
		#400 //152184900.0 * 1.4653913e+37 = 1.0385274e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111100011100010010100011110010;
		b = 32'b11111110000110001101011011010001;
		correct = 32'b00111101110010011111011110010011;
		#400 //-5.008696e+36 * -5.078951e+37 = 0.09861674
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111010100101100100100100011110;
		b = 32'b01100010000000101110011011100000;
		correct = 32'b01011000000100101111010000111101;
		#400 //3.9016376e+35 * 6.0367826e+20 = 646310800000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111000111011001001010110001;
		b = 32'b00110101111001000010111010010111;
		correct = 32'b01010000101100001100100001110001;
		#400 //40338.69 * 1.7000883e-06 = 23727410000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100010010101011110100010010010;
		b = 32'b11010011000000100100001110010000;
		correct = 32'b10001110110100100011000011011101;
		#400 //2.8990005e-18 * -559479260000.0 = -5.181605e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000101101000000010011111011;
		b = 32'b10001000011101101101001010011001;
		correct = 32'b01100111101110101011011010000011;
		#400 //-1.3098139e-09 * -7.427549e-34 = 1.7634538e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111101000110100011110011100101;
		b = 32'b11111010010000001010010100001011;
		correct = 32'b01000010010011001111011001010111;
		#400 //-1.2813581e+37 * -2.5006712e+35 = 51.240566
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110010000000000001001111100111;
		b = 32'b11001010000011001111010111000100;
		correct = 32'b11100111011010001001101010110001;
		#400 //2.536841e+30 * -2309489.0 = -1.0984426e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001111000001110101100101001110;
		b = 32'b11110101011111000100101111010111;
		correct = 32'b00011001000010010101010111110110;
		#400 //-2270776800.0 * -3.198235e+32 = 7.100094e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011010100111111100000100110110;
		b = 32'b10111000101000110100000010001100;
		correct = 32'b11100001011110101000010000000000;
		#400 //2.248348e+16 * -7.7844685e-05 = -2.8882485e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010001101010001100111001001001;
		b = 32'b00110110101010100110000011010000;
		correct = 32'b01011010011111011010001100110000;
		#400 //90626925000.0 * 5.0776653e-06 = 1.7848149e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010010110101001010111011001101;
		b = 32'b01010011001100010000011110001001;
		correct = 32'b10111111000110011100011101101001;
		#400 //-456732870000.0 * 760335600000.0 = -0.600699
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100100010001000101111111001000;
		b = 32'b00110010001010001001011101001100;
		correct = 32'b11110001100101010001100000001010;
		#400 //-1.4489854e+22 * 9.813288e-09 = -1.4765545e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100000111011111101111011101110;
		b = 32'b10111111101011001011111111111111;
		correct = 32'b00100000101100011011101111001001;
		#400 //-4.0635697e-19 * -1.3496093 = 3.0109232e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101111101100111001111110110000;
		b = 32'b10011010101011110000100110000000;
		correct = 32'b11010100100000110101101010100111;
		#400 //3.2673375e-10 * -7.239365e-23 = -4513293000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111011000100011001110000001000;
		b = 32'b01111010001000001000010001011101;
		correct = 32'b11000000011010000011100110001010;
		#400 //-7.560477e+35 * 2.0836304e+35 = -3.628512
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110100001000011011010101010001;
		b = 32'b00111100010011111000100010111010;
		correct = 32'b01110111010001110111100011101101;
		#400 //5.1247395e+31 * 0.0126668755 = 4.0457802e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101001100010101111001101010010;
		b = 32'b11011010011111101101100110001010;
		correct = 32'b10001110100010111001001111011110;
		#400 //6.1706404e-14 * -1.7933458e+16 = -3.4408536e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100111111111100000111000111110;
		b = 32'b11001001110010001001010000011010;
		correct = 32'b11011101101000100010000001101011;
		#400 //2.3994876e+24 * -1643139.2 = -1.4603069e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001001101010000101110011100001;
		b = 32'b10111001010110001110000001110011;
		correct = 32'b01001111110001101011110000000100;
		#400 //-1379228.1 * -0.00020682979 = 6668421000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000010110001000001110001010000;
		b = 32'b00100101110100100001011111000100;
		correct = 32'b11011100011011101111011001101000;
		#400 //-98.0553 * 3.6445297e-16 = -2.6904788e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100011101011110011010100011101;
		b = 32'b11101101001000111110001111000110;
		correct = 32'b10110110000010001101011011011100;
		#400 //6.464015e+21 * -3.1700886e+27 = -2.0390644e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100001101111011011101110110101;
		b = 32'b01011101010010011011000111100010;
		correct = 32'b11000011111100001101000101011010;
		#400 //-4.3749504e+20 * 9.083529e+17 = -481.63556
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010110111100101011010010001001;
		b = 32'b00000111111011110000010000001000;
		correct = 32'b01001110100000011111100111001111;
		#400 //3.9211142e-25 * 3.5963093e-34 = 1090316200.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101011111101100010011011100111;
		b = 32'b01001010001001010000000001001111;
		correct = 32'b11100001001111101111001111101110;
		#400 //-5.9515893e+26 * 2703379.8 = -2.2015365e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101101011101011100100110001001;
		b = 32'b11111111110100011100010011101000;
		correct = 32'b11111111110100011100010011101000;
		#400 //-4.7542168e+27 * nan = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010111010110100100111101101011;
		b = 32'b01011011111001010010100010100000;
		correct = 32'b00111010111100111110000110000000;
		#400 //240034630000000.0 * 1.29004875e+17 = 0.0018606633
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100010000010001100100110100000;
		b = 32'b11110110000110001000110010000000;
		correct = 32'b10101011011001011000110011011111;
		#400 //6.3082145e+20 * -7.7351445e+32 = -8.155264e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000001111000100101111011011000;
		b = 32'b11000001100110110101101101001110;
		correct = 32'b00111111101110101000001001010001;
		#400 //-28.29631 * -19.419582 = 1.457102
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100101111000101010110011111111;
		b = 32'b11001011101100000110100011111011;
		correct = 32'b01011001101001000111100011001101;
		#400 //-1.33805755e+23 * -23122422.0 = 5786840000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011010110111010000111010101100;
		b = 32'b10111111001101000110100001010011;
		correct = 32'b11011011000111001101011101011011;
		#400 //3.111105e+16 * -0.70471686 = -4.4146882e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101000001100011001010011010001;
		b = 32'b01001101011000100110011001100011;
		correct = 32'b10011010010010001100110001111000;
		#400 //-9.857743e-15 * 237397550.0 = -4.15242e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000011110000011000111100000010;
		b = 32'b11000000110010101000101100111101;
		correct = 32'b01000010011101001010010010101111;
		#400 //-387.11725 * -6.329497 = 61.160824
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101111001001111011101101010011;
		b = 32'b00111101100110101110000111110001;
		correct = 32'b00110001000010101001111001110100;
		#400 //1.5255112e-10 * 0.07562626 = 2.0171713e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100101111000010111100010010100;
		b = 32'b01000110001001010001001100110001;
		correct = 32'b11011111001011101101010011010111;
		#400 //-1.3309459e+23 * 10564.798 = -1.259793e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000110010010101000101001001010;
		b = 32'b00100110100100111001111000101001;
		correct = 32'b00011111001011111001111110011000;
		#400 //3.8093576e-35 * 1.0243043e-15 = 3.7189704e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100110101010010110000101000011;
		b = 32'b01100001101100011100011100001100;
		correct = 32'b01000100011100111110100001001110;
		#400 //3.9993705e+23 * 4.0992707e+20 = 975.62976
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001001101010001101001000101001;
		b = 32'b10100110001110000111100001110000;
		correct = 32'b01100010111010100100100001000100;
		#400 //-1382981.1 * -6.4001047e-16 = 2.1608727e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101011111111001110010011100011;
		b = 32'b01000100100110100001100011110001;
		correct = 32'b01100110110100100001000010010110;
		#400 //6.114604e+26 * 1232.7794 = 4.9600146e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010011010010101011010000000000;
		b = 32'b10111001101011001001011110011101;
		correct = 32'b10011001000101100101010011001010;
		#400 //2.5584731e-27 * -0.00032919357 = -7.771941e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101101000000110010100100011011;
		b = 32'b00110110000010011101001111101011;
		correct = 32'b10110110011100111001110111001001;
		#400 //-7.455615e-12 * 2.0537943e-06 = -3.6301665e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010101001010101111101010110101;
		b = 32'b11001011001000001001001010001101;
		correct = 32'b00001001100010000100101110111010;
		#400 //-3.4529e-26 * -10523277.0 = 3.2812022e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011010010010111001101011000011;
		b = 32'b00111010011101101100000011110011;
		correct = 32'b01011111010100110011101111100100;
		#400 //1.4327396e+16 * 0.0009412907 = 1.522101e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111001011011111101000101000000;
		b = 32'b01111001011100110011000101011000;
		correct = 32'b10111111011111000111001001100111;
		#400 //-7.782519e+34 * 7.892056e+34 = -0.98612064
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001111001011001001010111100111;
		b = 32'b10111000011111111011111000001110;
		correct = 32'b01010110001011001100001001101000;
		#400 //-2895505200.0 * -6.097374e-05 = 47487742000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010001000010000101110010001111;
		b = 32'b01101010011110000101010111100101;
		correct = 32'b00100110000011001001000111110100;
		#400 //36604277000.0 * 7.5054807e+25 = 4.877006e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101101011111100000001000110110;
		b = 32'b10000101001000101111111010010101;
		correct = 32'b01100111110001110111100101000011;
		#400 //-1.4438719e-11 * -7.663963e-36 = 1.8839756e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101001101101011001111000110111;
		b = 32'b10011010111000101000111101101010;
		correct = 32'b11001110010011010011011111001001;
		#400 //8.0654606e-14 * -9.370311e-23 = -860746300.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011000101101000011001011101000;
		b = 32'b00100110011101000101110001011111;
		correct = 32'b10110001101111001100100000101100;
		#400 //-4.658031e-24 * 8.477969e-16 = -5.494277e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010001110001010001110101111010;
		b = 32'b11001010000110111000010011111010;
		correct = 32'b00000111001000100011110000111011;
		#400 //-3.1099286e-28 * -2548030.5 = 1.2205226e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001010010110001001101011001101;
		b = 32'b01101011111101111010100011101100;
		correct = 32'b00011101110111111110011000100111;
		#400 //3548851.2 * 5.9880478e+26 = 5.926558e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001110010010101110010101101110;
		b = 32'b11010101110011111100010000011000;
		correct = 32'b00110111111110011111111111101011;
		#400 //-851008400.0 * -28555140000000.0 = 2.9802284e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000100000111001101100110011000;
		b = 32'b10001001011000111110101010101100;
		correct = 32'b10111010001100000010110100111000;
		#400 //1.8437626e-36 * -2.7434473e-33 = -0.00067206053
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100100001010100000001101101100;
		b = 32'b11111110110010101000101111100100;
		correct = 32'b00100100110101101110000110010110;
		#400 //-1.2544772e+22 * -1.346152e+38 = 9.3189863e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100110100011101000001111001010;
		b = 32'b11010011001001110001110000111111;
		correct = 32'b01010010110110100101001001010010;
		#400 //-3.3650356e+23 * -717733400000.0 = 468842000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101110010101011100111100011110;
		b = 32'b11011011110001110111001100000100;
		correct = 32'b01010010000010010011011100110100;
		#400 //-1.6542674e+28 * -1.1227996e+17 = 147334170000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110100001001010110011101010100;
		b = 32'b11010001110101010111111000101001;
		correct = 32'b11100001110001100101011000001001;
		#400 //5.24185e+31 * -114618080000.0 = -4.5733185e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010110000001110001000100100000;
		b = 32'b01010011000100111111100010101101;
		correct = 32'b00000010011010011010110010100101;
		#400 //1.0910617e-25 * 635532300000.0 = 1.7167683e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000001101011000011001010101110;
		b = 32'b11111101111101000001001001110101;
		correct = 32'b10000011001101001001110100000101;
		#400 //21.524746 * -4.0553433e+37 = -5.3077495e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110010011011000010010011010100;
		b = 32'b00100010111100011000100011111010;
		correct = 32'b11001110111110100100100100110011;
		#400 //-1.3745382e-08 * 6.546821e-18 = -2099550600.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011010101000011100100101001111;
		b = 32'b01011101110100000111001101000010;
		correct = 32'b10111100010001101011000100001101;
		#400 //-2.2769406e+16 * 1.8775527e+18 = -0.012127173
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001111010000100111011101010000;
		b = 32'b00101010110100010000100111000010;
		correct = 32'b01100011111011100010011101111100;
		#400 //3262599200.0 * 3.713263e-13 = 8.7863405e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100011110111111111011001001010;
		b = 32'b01111011010000100101100001111100;
		correct = 32'b10101000000100111000000110001000;
		#400 //-8.262742e+21 * 1.0091003e+36 = -8.188227e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100101110010111000110011010011;
		b = 32'b11001000100100000110001010011101;
		correct = 32'b00011100101101000111001101100001;
		#400 //-3.5310313e-16 * -295700.9 = 1.1941226e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100011100001001010110100100010;
		b = 32'b01010101110001101110110100001011;
		correct = 32'b10001101001010101011111000011011;
		#400 //-1.4384793e-17 * 27340174000000.0 = -5.2614126e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110101100101010010010000110011;
		b = 32'b01101011110100100001111000101110;
		correct = 32'b01001001001101011011010101011110;
		#400 //3.7811838e+32 * 5.080339e+26 = 744277.9
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101101000000100111110000011011;
		b = 32'b10110000101010110010101011000110;
		correct = 32'b00111011110000110010011110101011;
		#400 //-7.417201e-12 * -1.2454044e-09 = 0.0059556565
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001000110111101101110001101010;
		b = 32'b00110011100010101111111010110001;
		correct = 32'b01010100110011010011101101101000;
		#400 //456419.3 * 6.472454e-08 = 7051719700000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111101001011111010000100110010;
		b = 32'b10001100110110100110100110100000;
		correct = 32'b11101111110011011101101010111010;
		#400 //0.042878337 * -3.365179e-31 = -1.274177e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011001001000110110111101011110;
		b = 32'b10000100111000000110000000100011;
		correct = 32'b11010011101110100111100001100100;
		#400 //8.449393e-24 * -5.2750435e-36 = -1601767500000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110100101010111111000010010001;
		b = 32'b11011011010110111111110101000100;
		correct = 32'b00011000110010000001010111000100;
		#400 //-3.2026267e-07 * -6.192149e+16 = 5.1720766e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001010110001010111011011111100;
		b = 32'b00010111011000011101001010101001;
		correct = 32'b00110010110111111101101000110011;
		#400 //1.9015167e-32 * 7.296731e-25 = 2.6059842e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001000001011001001011011001111;
		b = 32'b10111010101010011111010001001101;
		correct = 32'b00001101000000011111110000000000;
		#400 //-5.193664e-34 * -0.0012966484 = 4.005453e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101011011111100100000010101001;
		b = 32'b10101001111000000111001011100101;
		correct = 32'b01000001000100001111111100100110;
		#400 //-9.032866e-13 * -9.967529e-14 = 9.062292
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011010111110100000001001101100;
		b = 32'b01010001100100001010101011101110;
		correct = 32'b01001000110111010011010001111000;
		#400 //3.5185704e+16 * 77667880000.0 = 453027.75
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000010110011111011010011000010;
		b = 32'b10100110010011011011101110101001;
		correct = 32'b11011100000000010011101001000001;
		#400 //103.85304 * -7.137799e-16 = -1.4549729e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111001000110011111010110111000;
		b = 32'b10001100100010010111011110110010;
		correct = 32'b01101100000011110101101100111111;
		#400 //-0.00014682754 * -2.1180231e-31 = 6.9322916e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010010110011100001101101000011;
		b = 32'b00011000111001001011010101000011;
		correct = 32'b00111001011001101011001110001101;
		#400 //1.3007148e-27 * 5.9119646e-24 = 0.00022001397
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000010011101110011010100011101;
		b = 32'b01010100011011001111101110100101;
		correct = 32'b10101101100001011000010111000001;
		#400 //-61.80187 * 4071336700000.0 = -1.5179748e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000001000101101111111111101011;
		b = 32'b00001001101111110111100110001111;
		correct = 32'b11110110110010011110001010010110;
		#400 //-9.43748 * 4.609589e-33 = -2.0473582e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111111010100001011011111100110;
		b = 32'b01100010111100101011101011011100;
		correct = 32'b10011011110111000010000100000111;
		#400 //-0.81530607 * 2.2387884e+21 = -3.641729e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011001000111010101010101101;
		b = 32'b10001100001000010000110001101010;
		correct = 32'b01111110100000100001010010111000;
		#400 //-10726061.0 * -1.2406725e-31 = 8.645361e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101001110011001000100011010111;
		b = 32'b11100100001000111010010101111010;
		correct = 32'b10000101000111111111101101001101;
		#400 //9.083158e-14 * -1.2074973e+22 = -7.522301e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011011111011110111110000010011;
		b = 32'b10101100011101001011010001100111;
		correct = 32'b01101110111110101000100111111101;
		#400 //-1.3481788e+17 * -3.477463e-12 = 3.8769035e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011110010010100101000100011010;
		b = 32'b01011001110100110010011110111010;
		correct = 32'b01000011111101010100100011011000;
		#400 //3.6446155e+18 * 7429362500000000.0 = 490.5691
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001011101110000111010101110111;
		b = 32'b00010010100010011011011111101011;
		correct = 32'b00111000101010110111000100101011;
		#400 //7.1050963e-32 * 8.691255e-28 = 8.1749946e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111110010010111010100110011111;
		b = 32'b11010000011000010110100111111111;
		correct = 32'b01101101011001110100110000010000;
		#400 //-6.76785e+37 * -15127281000.0 = 4.473937e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000010111000010101111010001000;
		b = 32'b00100110101100111011000000011101;
		correct = 32'b10011011101000001000101001111001;
		#400 //-3.3115037e-37 * 1.2468356e-15 = -2.6559265e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011000010000111101110011001000;
		b = 32'b00011111100111111110111111010000;
		correct = 32'b01111000000111001100000001111100;
		#400 //861412060000000.0 * 6.7735856e-20 = 1.2717224e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011111001001111010000010010101;
		b = 32'b01100110110101100110011100101001;
		correct = 32'b10110111110010000010011000110010;
		#400 //-1.2078818e+19 * 5.062447e+23 = -2.3859644e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001000011010001100010101010010;
		b = 32'b10111111110100110101010011010000;
		correct = 32'b10001000000011001111110001001101;
		#400 //7.004691e-34 * -1.6510258 = -4.2426296e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110101111001011001101011101101;
		b = 32'b01011000010011100001111000101010;
		correct = 32'b11011101000011101001010111110011;
		#400 //-5.821183e+32 * 906515800000000.0 = -6.421491e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100001110001101010010001111001;
		b = 32'b10101100000101101110011010101100;
		correct = 32'b01110101001010000111111011111111;
		#400 //-4.5803835e+20 * -2.144433e-12 = 2.1359416e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011110010011010110000000111100;
		b = 32'b10101101101101001001010000001010;
		correct = 32'b00110000000100011001001111010001;
		#400 //-1.08725104e-20 * -2.0529373e-11 = 5.296075e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011110111111110010010111101110;
		b = 32'b10110100011111011000010110110111;
		correct = 32'b10101010000000001101001000100100;
		#400 //2.7014863e-20 * -2.3611106e-07 = -1.1441591e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110011001100010010001011011111;
		b = 32'b01000100111101000001111101010010;
		correct = 32'b00101101101110011100000100110100;
		#400 //4.124274e-08 * 1952.9788 = 2.1117864e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100101100101111011000000000000;
		b = 32'b10101111101111100101001101011111;
		correct = 32'b11110101010011000000011101111100;
		#400 //8.95405e+22 * -3.4620037e-10 = -2.5863778e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100100111011000111000011111000;
		b = 32'b10101101110001100100011010011111;
		correct = 32'b11110110100110001010001101100110;
		#400 //3.4892575e+22 * -2.2541356e-11 = -1.547936e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111101001000110011111011111110;
		b = 32'b01010111101110010000110111001110;
		correct = 32'b11100100111000011101010011011001;
		#400 //-1.3561952e+37 * 406937900000000.0 = -3.3326838e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101011110111110100100001010010;
		b = 32'b10000111010001111001001100101011;
		correct = 32'b01100100000011110011010010001000;
		#400 //-1.5865176e-12 * -1.5014345e-34 = 1.0566679e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010000100010110111011101111001;
		b = 32'b01001101101001110101101010001101;
		correct = 32'b11000010010101010101011101100101;
		#400 //-18718902000.0 * 350966180.0 = -53.335346
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110110001001101011001011100110;
		b = 32'b01001001110110010010001011101001;
		correct = 32'b00101011110001001000100011110110;
		#400 //2.484006e-06 * 1778781.1 = 1.3964652e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000110011000111010001000101101;
		b = 32'b01111001101011011001100011010001;
		correct = 32'b00001100001001111101011111100100;
		#400 //14568.544 * 1.1267086e+35 = 1.2930179e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000001001010011101011101011110;
		b = 32'b10100101010100010100010011011000;
		correct = 32'b00011011010011111100010010010110;
		#400 //-3.1194916e-38 * -1.8151185e-16 = 1.7186159e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100010001101100111101000111000;
		b = 32'b10010011010101110101010001100100;
		correct = 32'b01001110010110001111000101011100;
		#400 //-2.4730301e-18 * -2.7178423e-27 = 909924100.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010111010101110100010110000001;
		b = 32'b10110001100101101010001100001001;
		correct = 32'b11100101001101101110101111110101;
		#400 //236693520000000.0 * -4.3841095e-09 = -5.398896e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001100110110100000001001100010;
		b = 32'b01110100110011001111110011111000;
		correct = 32'b00010111100010000010000101111001;
		#400 //114299660.0 * 1.2992668e+32 = 8.797244e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110000000101010100100001101000;
		b = 32'b11010110111100110001110000011001;
		correct = 32'b11011000100111010011001010111011;
		#400 //1.848032e+29 * -133651000000000.0 = -1382729700000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100000000110011101000001000110;
		b = 32'b01010000010110010001110000110001;
		correct = 32'b11001111001101010101110110001110;
		#400 //-4.4333743e+19 * 14570014000.0 = -3042807300.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011000010101111010111100100010;
		b = 32'b11101010011001110101011001010011;
		correct = 32'b10101101011011101010110110011010;
		#400 //948588760000000.0 * -6.991738e+25 = -1.3567281e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110101010111010110001111111101;
		b = 32'b00111011101001101010011001111101;
		correct = 32'b10111001001010100000101101101100;
		#400 //-8.247442e-07 * 0.005085765 = -0.00016216718
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101000010010110000010100001001;
		b = 32'b11010110111110000101100101000101;
		correct = 32'b11010000110100010100011001000001;
		#400 //3.834933e+24 * -136531150000000.0 = -28088338000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111011001000111100001000110;
		b = 32'b10110100100111011010100100110011;
		correct = 32'b11010010001110010111110011001111;
		#400 //58488.273 * -2.9366637e-07 = -199165720000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001001000100011101110111010000;
		b = 32'b11111011000110011100000101100100;
		correct = 32'b10001101011100101101110101110000;
		#400 //597469.0 * -7.9834385e+35 = -7.4838553e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100001011011010111100101101011;
		b = 32'b11011000011101101101111010111101;
		correct = 32'b10001000011101100100000110111001;
		#400 //8.045942e-19 * -1085746060000000.0 = -7.410519e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111000100101101110001110101;
		b = 32'b10110001110111011010110100011001;
		correct = 32'b01000100101010011001100111001111;
		#400 //-8.753607e-06 * -6.4516255e-09 = 1356.8065
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101000111001011000100001000011;
		b = 32'b11011100010111101101100101111001;
		correct = 32'b11001100000000111101011010100100;
		#400 //8.671484e+24 * -2.5090623e+17 = -34560656.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000101111011001110110110110001;
		b = 32'b11110010110100110110000101000010;
		correct = 32'b00010010100011110111100010000110;
		#400 //-7581.7114 * -8.373621e+30 = 9.05428e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100010101110110101111101010100;
		b = 32'b00011111000001001011101101101110;
		correct = 32'b01000011001101001011000100110100;
		#400 //5.0787384e-18 * 2.8107125e-20 = 180.6922
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000100011001011110001110001100;
		b = 32'b10110000010000000011101110111111;
		correct = 32'b00010011100110010001001010111011;
		#400 //-2.7023305e-36 * -6.99341e-10 = 3.86411e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110001000000111000101100101010;
		b = 32'b11011100000110011111011101011101;
		correct = 32'b00010100010110101011011111000011;
		#400 //-1.9142115e-09 * -1.733506e+17 = 1.1042428e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000010011100100101101011000001;
		b = 32'b10000111100100110110111000001111;
		correct = 32'b10111010010100100110101000010110;
		#400 //1.7805397e-37 * -2.2182788e-34 = -0.00080266723
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001001100001110010010100010010;
		b = 32'b11010001011110110011110111011011;
		correct = 32'b00110111100010011011010001010010;
		#400 //-1107106.2 * -67442160000.0 = 1.641564e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001000110101100110101111011001;
		b = 32'b01101101110001010000010111011101;
		correct = 32'b00011010100010110100110110011111;
		#400 //439134.78 * 7.6219544e+27 = 5.7614456e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000000000111101100111111111111;
		b = 32'b00101111010110010011100011011001;
		correct = 32'b11010000001110110010100111001110;
		#400 //-2.481445 * 1.9756231e-10 = -12560316000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010011010010010101111101111111;
		b = 32'b11110011110100010000110100101001;
		correct = 32'b10011110111101101001100011100100;
		#400 //864890600000.0 * -3.3125518e+31 = -2.6109497e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001001101100011101110111010000;
		b = 32'b00001100100011110001101110011100;
		correct = 32'b11111100100111110001011011010011;
		#400 //-1457082.0 * 2.2049255e-31 = -6.608305e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000101011010111001010010110110;
		b = 32'b00001100100111000111110111101001;
		correct = 32'b00111000010000001011000010001100;
		#400 //1.1076961e-35 * 2.4111385e-31 = 4.594079e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101000100001000001001001111000;
		b = 32'b01110011011011110010101100100100;
		correct = 32'b10110100100011010101110111100001;
		#400 //-4.9895445e+24 * 1.8948882e+31 = -2.6331602e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111101110110000111001100100;
		b = 32'b01101011101010101111111010101010;
		correct = 32'b00011011100011000000010111100001;
		#400 //95772.78 * 4.1344e+26 = 2.3164856e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101100100111011000101111000001;
		b = 32'b11100100010101110000111001011011;
		correct = 32'b01000111101110111000101001100111;
		#400 //-1.5236906e+27 * -1.5868338e+22 = 96020.805
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111110100000111011101011001010;
		b = 32'b01100101011111000010011000110110;
		correct = 32'b10011000100001011011110111001011;
		#400 //-0.25728446 * 7.4421326e+22 = -3.4571336e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010101101011100110010101001101;
		b = 32'b00111111101101010010010100101010;
		correct = 32'b11010101011101100111011000100001;
		#400 //-23968763000000.0 * 1.4151967 = -16936701000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111001000011000100010101001000;
		b = 32'b10100100010001111010011101010101;
		correct = 32'b01010100001100111101101110011110;
		#400 //-0.0001337725 * -4.3292982e-17 = 3089934800000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111011000001000110010100111010;
		b = 32'b01101110010001100001011111011010;
		correct = 32'b00001100001010110001100011101111;
		#400 //0.0020201937 * 1.5326717e+28 = 1.3180864e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101100100000111111000111110001;
		b = 32'b01010011110111110101101000000111;
		correct = 32'b11011000000101110011101101101011;
		#400 //-1.2760945e+27 * 1918576200000.0 = -665125800000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101110001010101101110001011110;
		b = 32'b11100111100000101010000111111000;
		correct = 32'b00000110001001110110101011011010;
		#400 //-3.884925e-11 * -1.2337909e+24 = 3.148771e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001010000111100011101000010000;
		b = 32'b00100000010011011001101110001110;
		correct = 32'b10101001010001010000000110110001;
		#400 //-7.6183436e-33 * 1.7415644e-19 = -4.3744254e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001111111100100111100101110011;
		b = 32'b00011001000000000000010011110110;
		correct = 32'b00110110011100100111000000001110;
		#400 //2.3909823e-29 * 6.618447e-24 = 3.6126035e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100111000101110101110001110010;
		b = 32'b00100010101100101000100000100100;
		correct = 32'b11000011110110010000101000011010;
		#400 //-2.1005574e-15 * 4.839114e-18 = -434.07892
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101111100011000111100010101011;
		b = 32'b01100100011001001001001010111100;
		correct = 32'b01001010100111010101001110100100;
		#400 //8.694756e+28 * 1.6865724e+22 = 5155282.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000101110110011100100111000001;
		b = 32'b00100010111010011011000101011110;
		correct = 32'b01100010011011101001001110111011;
		#400 //6969.219 * 6.334257e-18 = 1.10024255e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100101001100010111010001000001;
		b = 32'b01001000000001001100110011010000;
		correct = 32'b11011100101010110000101001000001;
		#400 //-5.237521e+22 * 135987.25 = -3.8514796e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010110010101010101011110101100;
		b = 32'b10000000000110101001100111011110;
		correct = 32'b01010110100000000101001000111110;
		#400 //-1.7233667e-25 * -2.44292e-39 = 70545360000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010011101010010111101110011111;
		b = 32'b11111101000001111100111111101101;
		correct = 32'b10010110000111111011101111011111;
		#400 //1455847000000.0 * -1.1282837e+37 = -1.2903199e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000011000110111010001001101100;
		b = 32'b10010111010111110111101000101100;
		correct = 32'b10101011001100100100100010110110;
		#400 //4.5736857e-37 * -7.220939e-25 = -6.333921e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101010101001100101011000111011;
		b = 32'b11111111110010001111100100000101;
		correct = 32'b11111111110010001111100100000101;
		#400 //-2.9547358e-13 * nan = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000011001010011101001010110010;
		b = 32'b11111100010001111111011010110011;
		correct = 32'b00000110010110010110100110111000;
		#400 //-169.82303 * -4.153083e+36 = 4.0890834e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000010011101110111110011110001;
		b = 32'b11001110011001001110111001001100;
		correct = 32'b00110011100010100110000000101111;
		#400 //-61.872013 * -960205600.0 = 6.4436215e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100101000000001000101110001001;
		b = 32'b10110000001000111111100100110011;
		correct = 32'b01110100010010001011000000101111;
		#400 //-3.7939805e+22 * -5.965319e-10 = 6.3600635e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110101001111011010101111111100;
		b = 32'b00100011011110100100001100001010;
		correct = 32'b01010001010000100000010101001101;
		#400 //7.0658257e-07 * 1.3566723e-17 = 52082037000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110000111001001011000000011101;
		b = 32'b11010111101100011111011011000100;
		correct = 32'b01011000101001000111101110101100;
		#400 //-5.6620392e+29 * -391346820000000.0 = 1446808600000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110110110000010010100010011001;
		b = 32'b01111100000011011010011001000110;
		correct = 32'b10111010001011101000101110101101;
		#400 //-1.9588608e+33 * 2.941945e+36 = -0.00066583866
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001001110100001010100001010110;
		b = 32'b11110100100001001001100010110100;
		correct = 32'b00010100110010010110110010100101;
		#400 //-1709322.8 * -8.404301e+31 = 2.0338666e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111011010011111010011010101100;
		b = 32'b11110000101010001101001010011001;
		correct = 32'b00001010000111010111000001111100;
		#400 //-0.0031685038 * -4.1798463e+29 = 7.580431e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011110011000001010110001110111;
		b = 32'b11111110100011111010111001100000;
		correct = 32'b10011111010010000010011100110100;
		#400 //4.0473614e+18 * -9.549251e+37 = -4.2384075e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111111110101010011100001000010;
		b = 32'b00111010110111011111101110110100;
		correct = 32'b01000100011101011110010011000101;
		#400 //1.6657794 * 0.0016935975 = 983.5745
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010001101100001000010100010000;
		b = 32'b01101111110000111001101111011001;
		correct = 32'b10100001011001110000010001111111;
		#400 //-94768330000.0 * 1.2107597e+29 = -7.8271795e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001100000111011000111001101000;
		b = 32'b00000001100001011111101010000011;
		correct = 32'b11001010000101101000011010001110;
		#400 //-1.2137694e-31 * 4.921595e-38 = -2466211.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100011101101111101010110001110;
		b = 32'b00010010100111110000100011100100;
		correct = 32'b01010000100100111111010111000010;
		#400 //1.9931344e-17 * 1.0036502e-27 = 19858854000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010011011010101001100001000011;
		b = 32'b11100101100111101000000110011100;
		correct = 32'b00101101001111010111000111000101;
		#400 //-1007576900000.0 * -9.35656e+22 = 1.0768668e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111001000111011001111110100011;
		b = 32'b00110111111011000011000110101100;
		correct = 32'b01000000101010101101011101001111;
		#400 //0.00015032156 * 2.8156523e-05 = 5.338783
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010011010110110110000111010111;
		b = 32'b00110011010011110110100110001001;
		correct = 32'b10011111100001110110001100010010;
		#400 //-2.7689925e-27 * 4.8291927e-08 = -5.733862e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110010101011101101110001000101;
		b = 32'b00100010101100000010110111111110;
		correct = 32'b11001111011111100001010101000101;
		#400 //-2.0356433e-08 * 4.775359e-18 = -4262806800.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101010101111110100011011011010;
		b = 32'b10000100001110001011001010000111;
		correct = 32'b11100110000001001000111101001000;
		#400 //3.397758e-13 * -2.1711072e-36 = -1.5649886e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100111000001101000101100111000;
		b = 32'b10111111110000010000111001111101;
		correct = 32'b01100110101100100110100011110011;
		#400 //-6.3536524e+23 * -1.5082546 = 4.212586e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111111100100100110011011110;
		b = 32'b01111111111100001110010110100000;
		correct = 32'b01111111111100001110010110100000;
		#400 //-2.8884442e-05 * nan = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010100010111010010000110100001;
		b = 32'b01101111000010010000100101011101;
		correct = 32'b10100100110011101000110010100010;
		#400 //-3799008000000.0 * 4.2410766e+28 = -8.95765e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010111100011101110000101010011;
		b = 32'b01011000011101000111110000101000;
		correct = 32'b00111110100101011001110000010101;
		#400 //314196820000000.0 * 1075256340000000.0 = 0.29220644
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110110011000011001101011000011;
		b = 32'b10111011111001000000101001000101;
		correct = 32'b11111001111111010100010000001011;
		#400 //1.1439509e+33 * -0.006959232 = -1.643789e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101001110010011011100011000111;
		b = 32'b01110011001011000110000101001001;
		correct = 32'b10110110000101011100100110100000;
		#400 //-3.0483335e+25 * 1.3657352e+31 = -2.2320091e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101111110101110110010110110011;
		b = 32'b01101010111100001010010011110000;
		correct = 32'b10000100011001010010010001010110;
		#400 //-3.9180534e-10 * 1.4546055e+26 = -2.6935505e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100011010000011000000100000001;
		b = 32'b00101101010001011110010111011111;
		correct = 32'b00110101011110100101000011100000;
		#400 //1.0489869e-17 * 1.1249195e-11 = 9.3249946e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000101000101100010000100010;
		b = 32'b11001001010000101110010100000110;
		correct = 32'b00100110110101011100110001011011;
		#400 //-1.1842796e-09 * -798288.4 = 1.4835235e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111000000011110110001000000101;
		b = 32'b11001110111101001001001100100100;
		correct = 32'b01101000100101100001010010111011;
		#400 //-1.1632602e+34 * -2051641900.0 = 5.669899e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111100110001011010100010010000;
		b = 32'b00110010011011001110010001110100;
		correct = 32'b01001001110101011001100111111010;
		#400 //0.024128228 * 1.3788952e-08 = 1749823.2
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011001011110001100111011000101;
		b = 32'b00100000011111111011000001000101;
		correct = 32'b01111000011110010001110001011011;
		#400 //4377071200000000.0 * 2.1657663e-19 = 2.0210266e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001010110101011100101001010101;
		b = 32'b10001100011011000001110000000001;
		correct = 32'b00111101111001111100110011111101;
		#400 //-2.0587263e-32 * -1.8189206e-31 = 0.11318395
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110000100101111100111100100011;
		b = 32'b10110100001111001110111111010011;
		correct = 32'b10111011110011011011000110011111;
		#400 //1.1045568e-09 * -1.7596112e-07 = -0.0062772776
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000010100001100001001101100110;
		b = 32'b10111011101000011000000110011110;
		correct = 32'b10000110010101001000010100111110;
		#400 //1.9700665e-37 * -0.0049287817 = -3.997066e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011110111000010001001010111000;
		b = 32'b10110110000101100110011010101001;
		correct = 32'b00101000001111111000110011100000;
		#400 //-2.3830544e-20 * -2.2411498e-06 = 1.0633177e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010101000011110001111101010;
		b = 32'b11101000000011000101010100101010;
		correct = 32'b00010010000100111010100111000001;
		#400 //-0.0012351249 * -2.6508092e+24 = 4.659426e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100100101110101010001011101011;
		b = 32'b11011110111011111000100111110111;
		correct = 32'b00000101010001110111011001000111;
		#400 //-8.0940635e-17 * -8.6302993e+18 = 9.378659e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011100010000101010110010100100;
		b = 32'b11000010011001110011111100100001;
		correct = 32'b01011001010101111000001101010010;
		#400 //-2.1918386e+17 * -57.81165 = 3791344300000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000010101101000000110011100101;
		b = 32'b11001110111100100010101111110110;
		correct = 32'b00110011001111100101010011011010;
		#400 //-90.025185 * -2031483600.0 = 4.4314994e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111101001010100111111101010111;
		b = 32'b11011010111111011101111001110011;
		correct = 32'b01100001101010111110110110111011;
		#400 //-1.4164372e+37 * -3.5728877e+16 = 3.9644044e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110101010100100001110000100110;
		b = 32'b11001011001000011100100110011011;
		correct = 32'b00101001101001100011101100011000;
		#400 //-7.827206e-07 * -10602907.0 = 7.382132e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010101000110000010100000101010;
		b = 32'b00101100111000000111101010001011;
		correct = 32'b10100111101011011000010111010101;
		#400 //-3.072784e-26 * 6.380068e-12 = -4.8162247e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001100100101111100000001000110;
		b = 32'b10111101010000000100001001011000;
		correct = 32'b11001110110010100000111111100001;
		#400 //79561260.0 * -0.04693827 = -1695019100.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010111110101100010010111011010;
		b = 32'b00101011111110001101011101000010;
		correct = 32'b10101011010111000100111100010011;
		#400 //-1.3838981e-24 * 1.7681206e-12 = -7.826944e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100110101000101001011100110110;
		b = 32'b01011001110011011011111101001011;
		correct = 32'b01001100010010100100110101111010;
		#400 //3.8390636e+23 * 7239087400000000.0 = 53032424.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100001101001111110100110001011;
		b = 32'b00101011111010101010101111101110;
		correct = 32'b11110101001101110010110001010101;
		#400 //-3.8717935e+20 * 1.667442e-12 = -2.3219958e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111100001110100100100010011011;
		b = 32'b00100110010010010110110110101100;
		correct = 32'b01010101011011001100000010001100;
		#400 //0.01136985 * 6.9884517e-16 = 16269483000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100110010101111101010010101010;
		b = 32'b11011110001101000000100001001001;
		correct = 32'b01000111100110010111001110111000;
		#400 //-2.5480794e+23 * -3.2431747e+18 = 78567.44
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110011111101100110000010001111;
		b = 32'b10010000010111111010001000010000;
		correct = 32'b11100011000011010000010010011010;
		#400 //1.14728316e-07 * -4.4103844e-29 = -2.6013225e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110000000101010001111110000010;
		b = 32'b01101101010101000110000100000000;
		correct = 32'b01000010001100111100000001111011;
		#400 //1.8460543e+29 * 4.1080055e+27 = 44.93797
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011111110000101001000101010100;
		b = 32'b00001110100000010101001010001111;
		correct = 32'b01010000110000001001001111110110;
		#400 //8.240262e-20 * 3.1880456e-30 = 25847378000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000011010110000010101000010111;
		b = 32'b10111100010111011110000000001001;
		correct = 32'b01000110011110010110100100110100;
		#400 //-216.16441 * -0.013542184 = 15962.301
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110100111011110000000111100100;
		b = 32'b11001000000100001010111010101111;
		correct = 32'b00101100010100110111001011110100;
		#400 //-4.4518595e-07 * -148154.73 = 3.0048715e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110111000100100000100101011101;
		b = 32'b11000111110100011110001101110001;
		correct = 32'b11101110101100100001111011000011;
		#400 //2.9619736e+33 * -107462.88 = -2.756276e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010111000000011011011001011100;
		b = 32'b11011000001111100100110111001101;
		correct = 32'b10111110001011100111110111000000;
		#400 //142620230000000.0 * -836965440000000.0 = -0.17040157
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010110000101001001000111110001;
		b = 32'b11100010010010110011100111000011;
		correct = 32'b00110011001110110010011010111100;
		#400 //-40838634000000.0 * -9.372128e+20 = 4.357456e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010110011001100001100100001011;
		b = 32'b01001001000100010111110110100010;
		correct = 32'b11001100110010100110111110001010;
		#400 //-63248810000000.0 * 595930.1 = -106134610.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111000100100110011100000111011;
		b = 32'b00111100011101100010101111100101;
		correct = 32'b10111011100110010001100011110100;
		#400 //-7.01998e-05 * 0.015025114 = -0.004672164
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110001101111111000011011110011;
		b = 32'b01000111011010111011111111101100;
		correct = 32'b10101001110011111111101010010110;
		#400 //-5.5741736e-09 * 60351.92 = -9.2361164e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110110111101100100011011101100;
		b = 32'b11101001111001100010010001100011;
		correct = 32'b01001100100010001111100101010000;
		#400 //-2.4975459e+33 * -3.4778096e+25 = 71813760.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101111010001111111000000111010;
		b = 32'b00001000000101110000101111111111;
		correct = 32'b11100110101010010110111001111110;
		#400 //-1.818429e-10 * 4.545401e-34 = -4.0005908e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010110100010001001111100001110;
		b = 32'b10101000000001110010001100001011;
		correct = 32'b11101110000000010110011111110001;
		#400 //75108360000000.0 * -7.501604e-15 = -1.0012306e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110000111111010011010001000001;
		b = 32'b01000001000011101110001111010011;
		correct = 32'b11101111011000101101000110011110;
		#400 //-6.2690303e+29 * 8.930621 = -7.0197024e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001101110111100110011111010101;
		b = 32'b00011011000110001110111000001011;
		correct = 32'b11110010001110100010011001110000;
		#400 //-466418340.0 * 1.2650061e-22 = -3.6870835e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000011001011101110000000101;
		b = 32'b10100100110111011111011101100000;
		correct = 32'b01001011000001001000110100111100;
		#400 //-8.362238e-10 * -9.626254e-17 = 8686908.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101010101111001010101111101010;
		b = 32'b00111000101100001011010001110000;
		correct = 32'b10110001100010001010101100011001;
		#400 //-3.3514798e-13 * 8.425943e-05 = -3.9775725e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000110011000100100110101001001;
		b = 32'b00001101111000110010111111110011;
		correct = 32'b11110111111111110000000010010111;
		#400 //-14483.321 * 1.40014985e-30 = -1.03441224e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110110011101111000110110101110;
		b = 32'b01000110111111111010101100010111;
		correct = 32'b01101110111101111101111111100101;
		#400 //1.25524505e+33 * 32725.545 = 3.8356735e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101100110100010101000101111111;
		b = 32'b10100110101010011011010101110010;
		correct = 32'b01000101100111011101111111110111;
		#400 //-5.949185e-12 * -1.1775912e-15 = 5051.9956
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101000110101001110011110010101;
		b = 32'b10011001100110010101111010011110;
		correct = 32'b11001110101100011010111111100010;
		#400 //2.363716e-14 * -1.5858045e-23 = -1490547000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000110101011100101010011001100;
		b = 32'b00001100010101101001101001101100;
		correct = 32'b01111001110011111111010110101000;
		#400 //22314.398 * 1.653243e-31 = 1.3497349e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011000101010011101000110010101;
		b = 32'b10110111000111100011110100001010;
		correct = 32'b10100001000010010101111000001001;
		#400 //4.38971e-24 * -9.431746e-06 = -4.654186e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101111010011000111111100010011;
		b = 32'b10010101000010110110100011111001;
		correct = 32'b01011001101110111100001001100011;
		#400 //-1.8598838e-10 * -2.8153635e-26 = 6606194000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100111110001111100101100101111;
		b = 32'b01010101010110010011100100111100;
		correct = 32'b01010001111010110111010101101111;
		#400 //1.886998e+24 * 14927490000000.0 = 126410940000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110100010101101000101111111001;
		b = 32'b01111110011001010000000010001101;
		correct = 32'b00110101011011111101011100100110;
		#400 //6.7992585e+31 * 7.609902e+37 = 8.934752e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101010000011101111000001011011;
		b = 32'b10000101100101110000100000001110;
		correct = 32'b01100011111100100100100001110010;
		#400 //-1.2695524e-13 * -1.420293e-35 = 8.9386646e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000101110100100011010110000100;
		b = 32'b10111001111000110100000011000010;
		correct = 32'b00001011011011001100110011010001;
		#400 //-1.9767964e-35 * -0.00043345062 = 4.5606033e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010111001110100100110001101001;
		b = 32'b10101011010010000000110110101011;
		correct = 32'b00101011011011100110010111111110;
		#400 //-6.0196285e-25 * -7.107324e-13 = 8.469613e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100101011101101111011010111010;
		b = 32'b00101011110101001000100100010011;
		correct = 32'b00111001000101001011110000001011;
		#400 //2.1420693e-16 * 1.5101552e-12 = 0.00014184431
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100011100001001010100111111001;
		b = 32'b01111000000011010101000000101010;
		correct = 32'b00101010111100000101010011010001;
		#400 //4.894436e+21 * 1.1464684e+34 = 4.2691417e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000000110010100100011101011011;
		b = 32'b11111011101100111111001000011101;
		correct = 32'b00000100100011111110001011010010;
		#400 //-6.3212104 * -1.8686636e+36 = 3.382744e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011001010000101100111111001001;
		b = 32'b10110110110101110111100010010010;
		correct = 32'b11100001111001110111010001101100;
		#400 //3427163000000000.0 * -6.4215355e-06 = -5.3369837e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000011000101101110011010001100;
		b = 32'b01011111011111011110001111010001;
		correct = 32'b10100011000110000010011110011011;
		#400 //-150.90057 * 1.8294696e+19 = -8.248323e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100111000101001011101001000010;
		b = 32'b11101010100011101011011101000000;
		correct = 32'b10111100000001010110010001010001;
		#400 //7.023461e+23 * -8.626642e+25 = -0.008141593
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111100110101101111100111100000;
		b = 32'b00000011010001000000111101010000;
		correct = 32'b01111001000011000101100110000110;
		#400 //0.026242197 * 5.76168e-37 = 4.554608e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101101110010101000001001111010;
		b = 32'b11101111101001111110000001111100;
		correct = 32'b00111101100110100110011111111111;
		#400 //-7.8342136e+27 * -1.0391076e+29 = 0.07539367
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100000101111110110110111010101;
		b = 32'b10010100100111011010010010010100;
		correct = 32'b01001011100110110110111011011101;
		#400 //-3.242934e-19 * -1.5917863e-26 = 20372922.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010010001100111101011001101111;
		b = 32'b01110011011111111111010101101000;
		correct = 32'b10011110001100111101110111100000;
		#400 //-193099190000.0 * 2.0279131e+31 = -9.522064e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010100010110101011111100101000;
		b = 32'b11110100010001001100100000001001;
		correct = 32'b00011111100011100100100110101001;
		#400 //-3758039800000.0 * -6.236251e+31 = 6.02612e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000000100101110001101011101111;
		b = 32'b01100101011100101111010101000100;
		correct = 32'b10011010100111110011011101101101;
		#400 //-4.722038 * 7.1708565e+22 = -6.5850404e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010010011110101000001001110111;
		b = 32'b01000010010011110001110110101110;
		correct = 32'b01001111100110101101000101011011;
		#400 //268982670000.0 * 51.778984 = 5194823000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001100111101011101101011100110;
		b = 32'b01101101001000011100101010001001;
		correct = 32'b10011111010000101000000110110001;
		#400 //-128898860.0 * 3.129496e+27 = -4.1188376e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000000001100100110010101000010;
		b = 32'b11111010111111000000001011010011;
		correct = 32'b10000100101101010011100000100011;
		#400 //2.7874303 * -6.5425805e+35 = -4.260445e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110001011100100101011000101100;
		b = 32'b11100111101010000111111110111100;
		correct = 32'b01001001001110000001011100110110;
		#400 //-1.1999928e+30 * -1.5914277e+24 = 754035.4
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010101111010001110010110010;
		b = 32'b10110110110111000001101000010110;
		correct = 32'b01000011010110111111010010110001;
		#400 //-0.0014428108 * -6.5595477e-06 = 219.95583
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110010010111101001110111011011;
		b = 32'b01011101101100101100111101000110;
		correct = 32'b11010100000111110101101111100111;
		#400 //-4.4093765e+30 * 1.6105743e+18 = -2737766700000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100111111011100011110101100001;
		b = 32'b10101110111100111011100000001101;
		correct = 32'b00111000011110100011111010100110;
		#400 //-6.6124817e-15 * -1.10830546e-10 = 5.966299e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010101100000101001011100001100;
		b = 32'b11010001111110100011111001100000;
		correct = 32'b00000011000001011001100000001111;
		#400 //-5.274489e-26 * -134348540000.0 = 3.925974e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111111110010111100101111101010;
		b = 32'b00100001000110101111000000000001;
		correct = 32'b11011110001010000101110101000111;
		#400 //-1.5921605 * 5.249487e-19 = -3.0329828e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001000111111010000001100010011;
		b = 32'b01101111010111000101101010001111;
		correct = 32'b10011001000100101111100001111110;
		#400 //-518168.6 * 6.819618e+28 = -7.598206e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101010000111000100111010110011;
		b = 32'b00101000111001111110000110010011;
		correct = 32'b11000000101011001001000011001000;
		#400 //-1.3882888e-13 * 2.5743979e-14 = -5.3926735
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101110111100010111100001000011;
		b = 32'b11011011111000011001101010010001;
		correct = 32'b00010010100010010000000001111000;
		#400 //-1.0980774e-10 * -1.27003635e+17 = 8.646031e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011111010110110101110000000110;
		b = 32'b01111100110010111010011011001101;
		correct = 32'b00100010000010011101111101110000;
		#400 //1.5806515e+19 * 8.459355e+36 = 1.868525e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111111110101100000001110101010;
		b = 32'b10111100111011000001110100111101;
		correct = 32'b01000010011010000000100111110000;
		#400 //-1.6719868 * -0.028822536 = 58.009705
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100000110000000110110010010011;
		b = 32'b10110011111000011111111111001111;
		correct = 32'b01101100010110011111011111000110;
		#400 //-1.1092495e+20 * -1.052391e-07 = 1.0540279e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011001010111110011110010011110;
		b = 32'b00111001001010011100000011100000;
		correct = 32'b00011111101010000101010000001101;
		#400 //1.1541071e-23 * 0.00016188947 = 7.128982e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000111110101100011110100010111;
		b = 32'b10101110110101011101111000011001;
		correct = 32'b10011000100000000011100011011010;
		#400 //3.2235047e-34 * -9.725571e-11 = -3.314463e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111010000000001010000001011011;
		b = 32'b01101111100011000110001110110100;
		correct = 32'b11001001111010101000110011010000;
		#400 //-1.669666e+35 * 8.689687e+28 = -1921434.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000000110110011011101010001000;
		b = 32'b01100111111010100101111000010011;
		correct = 32'b10011000011011011101001101001011;
		#400 //-6.80402 * 2.2135382e+24 = -3.0738208e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010111011010001110000000100011;
		b = 32'b00011100111101111100101100111101;
		correct = 32'b11111001111100001001011001101100;
		#400 //-256049360000000.0 * 1.6397625e-21 = -1.5615027e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111010010100010100111101101110;
		b = 32'b01000010111001101010100110001111;
		correct = 32'b01110110111010000100110101101110;
		#400 //2.7170027e+35 * 115.33117 = 2.3558268e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101110100111111011111001000010;
		b = 32'b01000011000011000001011101110110;
		correct = 32'b01101011000100011111010010010100;
		#400 //2.4719062e+28 * 140.09164 = 1.7644923e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000000111100100111011100110011;
		b = 32'b11110010110010100111110100011000;
		correct = 32'b00001101100110010100010101010100;
		#400 //-7.5770507 * -8.021402e+30 = 9.446043e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001110011100000110101001000110;
		b = 32'b01010111001011011001110011000010;
		correct = 32'b00110110101100010100000010000100;
		#400 //1008374140.0 * 190888780000000.0 = 5.2825217e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111011010011101101000010110111;
		b = 32'b11011011001110011010011010001010;
		correct = 32'b01011111100011101001011110101000;
		#400 //-1.0738464e+36 * -5.2255982e+16 = 2.0549732e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101100000001010110001000111010;
		b = 32'b10011001001100010010101101111101;
		correct = 32'b01010010010000001011101101001000;
		#400 //-1.8954963e-12 * -9.159468e-24 = 206943940000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110111011010111110010101000011;
		b = 32'b01010000010101110101100111111010;
		correct = 32'b01100110100011000011011000000000;
		#400 //4.7845302e+33 * 14451993000.0 = 3.310637e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111011011001110111001001111000;
		b = 32'b00010010101111111111010110100100;
		correct = 32'b11101000000110100101010010100100;
		#400 //-0.0035316031 * 1.211435e-27 = -2.915223e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011000101100010011001001000001;
		b = 32'b10111101101000010001010001011000;
		correct = 32'b10011010100011001100111010011100;
		#400 //4.580417e-24 * -0.078652084 = -5.823644e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011101110111101011101001001010;
		b = 32'b10111001100000010000100001011001;
		correct = 32'b10100011110111001111000111111101;
		#400 //5.895553e-21 * -0.00024611017 = -2.3954934e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011000010101101000010011111011;
		b = 32'b11001110101001011110001100010111;
		correct = 32'b00001001001001011000011001110011;
		#400 //-2.772599e-24 * -1391561600.0 = 1.992437e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110100011101001110001000110001;
		b = 32'b01101010010111111110000100000111;
		correct = 32'b10001001100011000000001001010011;
		#400 //-2.2806559e-07 * 6.766328e+25 = -3.370596e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100110110101111111100101010101;
		b = 32'b00110011011110000000010101001100;
		correct = 32'b00110010110111101110110000011001;
		#400 //1.4986203e-15 * 5.7746817e-08 = 2.5951566e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011000011111100010010100100101;
		b = 32'b00011001000101110100110011010101;
		correct = 32'b11111110110101110000000111000101;
		#400 //-1117741950000000.0 * 7.822033e-24 = -1.428966e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010010100111101111010001101010;
		b = 32'b01001110010000000000001011111100;
		correct = 32'b10000011110100111110110101000010;
		#400 //-1.0031455e-27 * 805355260.0 = -1.2455937e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001101010100101001011000100010;
		b = 32'b01010110011001000011100011100100;
		correct = 32'b00110110011011000011011110111100;
		#400 //220815900.0 * 62733250000000.0 = 3.5199182e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111111100001010110011101010001;
		b = 32'b01011000000100001001100101010100;
		correct = 32'b00100110111011000010110111111001;
		#400 //1.0422155 * 635952850000000.0 = 1.638825e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100001110101010111101101010011;
		b = 32'b01010110000110101101111110110000;
		correct = 32'b00001011001100000111000000110011;
		#400 //1.4466085e-18 * 42571380000000.0 = 3.3980776e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001101001100001111011000101101;
		b = 32'b01001100000011010100001111010111;
		correct = 32'b00000000101000000101100000111011;
		#400 //5.453051e-31 * 37031772.0 = 1.472533e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101101010100101011101010100111;
		b = 32'b11100101000000001001010100100110;
		correct = 32'b11000111110100011100011000111000;
		#400 //4.0760938e+27 * -3.795089e+22 = -107404.44
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101100100010100011100100110000;
		b = 32'b10000110101110100111100101011100;
		correct = 32'b11100101001111011100001001100010;
		#400 //3.928545e-12 * -7.0143745e-35 = -5.600706e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101111001101000011100110101110;
		b = 32'b01011110011111101000110010010000;
		correct = 32'b00010000001101010100000010101010;
		#400 //1.6391397e-10 * 4.5855484e+18 = 3.574577e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111000001111011101100011000101;
		b = 32'b10000110001001100110010001111111;
		correct = 32'b11110001100100100000101011100001;
		#400 //4.5262994e-05 * -3.1294963e-35 = -1.4463348e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111101110100100000111010110001;
		b = 32'b10111101110001001111010100000000;
		correct = 32'b00111111100010001000001110000110;
		#400 //-0.102567084 * -0.096170425 = 1.0665138
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010000000001010010000010111110;
		b = 32'b01110010000111100110011000101101;
		correct = 32'b10011101010101110010100001001011;
		#400 //-8934062000.0 * 3.137418e+30 = -2.8475844e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111010100001000010011000011110;
		b = 32'b11001100101010010101100010010110;
		correct = 32'b11101101010001111100010011101000;
		#400 //3.4307815e+35 * -88786100.0 = -3.8640976e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001111001000001001111000101111;
		b = 32'b00100111000010000000100010110110;
		correct = 32'b11100111100101110010000111001001;
		#400 //-2694721300.0 * 1.8878514e-15 = -1.4274011e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111001000010111110000111100010;
		b = 32'b11011101011011011111111111000110;
		correct = 32'b11011011000101100111011001010110;
		#400 //4.539442e+34 * -1.0718527e+18 = -4.235136e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001110110010100011001110011000;
		b = 32'b11100011011011101010010011010101;
		correct = 32'b10101010110110001110100001000011;
		#400 //1696189400.0 * -4.4022025e+21 = -3.8530472e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001111110000111111100000001010;
		b = 32'b10011000011010100010110110101001;
		correct = 32'b00110110110101100011101011100100;
		#400 //-1.9324026e-29 * -3.0266844e-24 = 6.3845528e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011111110100010000011010100101;
		b = 32'b01010011010111010100010011001100;
		correct = 32'b01001011111100011101010111100110;
		#400 //3.0123815e+19 * 950342000000.0 = 31697868.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111001010001001101110000101011;
		b = 32'b00011100110001001110110000111100;
		correct = 32'b11011011111111111110101100011101;
		#400 //-0.00018774036 * 1.3031257e-21 = -1.4406926e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100110100011100000100110100001;
		b = 32'b10110100010100000100101000011001;
		correct = 32'b00110001101011101001001010010110;
		#400 //-9.855839e-16 * -1.9398466e-07 = 5.0807314e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010001100010011001001011001100;
		b = 32'b11101010100010000010000000011011;
		correct = 32'b10100110100000010101110010010001;
		#400 //73859170000.0 * -8.228276e+25 = -8.976263e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111001110111101110010101001101;
		b = 32'b10111000001111001110111011000110;
		correct = 32'b11000001000101110000001001110100;
		#400 //0.00042513982 * -4.5045068e-05 = -9.438099
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100000010011010101101110001000;
		b = 32'b00110011100101000000110100011110;
		correct = 32'b00101100001100011000101110001001;
		#400 //1.739446e-19 * 6.894173e-08 = 2.523067e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001111100100110000001010011001;
		b = 32'b11100010010010011111001011101101;
		correct = 32'b00101100101110100101101101100101;
		#400 //-4932842000.0 * -9.3132505e+20 = 5.296585e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011010111110100110110110110111;
		b = 32'b11000100100110001010010001001110;
		correct = 32'b11010101110100100000000000100001;
		#400 //3.5244688e+16 * -1221.1345 = -28862250000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011001101100010111000111000000;
		b = 32'b11000111100001000000101010011000;
		correct = 32'b10010001101011000000001101101000;
		#400 //1.8347314e-23 * -67605.19 = -2.7138914e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011011010011010010110010100001;
		b = 32'b01000101111111001100110011101000;
		correct = 32'b10010100110011111100010101101001;
		#400 //-1.6971623e-22 * 8089.6133 = -2.0979523e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001111011110111000110110111101;
		b = 32'b10101000110101000011100000010110;
		correct = 32'b10100110000101111011100110000011;
		#400 //1.2402553e-29 * -2.3561052e-14 = -5.2640064e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111101110101000101101110101001;
		b = 32'b00001001001010111010101101010100;
		correct = 32'b11110100000111100101011010100000;
		#400 //-0.10369045 * 2.0663934e-33 = -5.0179435e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101111101000001100111001111101;
		b = 32'b01000000111011001100010001011111;
		correct = 32'b01101110001011011101111010000000;
		#400 //9.953446e+28 * 7.398971 = 1.3452473e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000110101110110001010000111110;
		b = 32'b00010100001010111001111111101111;
		correct = 32'b10110010000010111000011010101011;
		#400 //-7.0371325e-35 * 8.664835e-27 = -8.121485e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010001001001111001110001111011;
		b = 32'b00011110010010001001100101001000;
		correct = 32'b00110010010101011110011011101011;
		#400 //1.3222196e-28 * 1.061961e-20 = 1.2450736e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000101101110111000001101000100;
		b = 32'b11111001101001110110100101001110;
		correct = 32'b10001011100011110101111010000101;
		#400 //6000.408 * -1.0865618e+35 = -5.5223814e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011111111001001011011111110010;
		b = 32'b00101001000101000101111101001010;
		correct = 32'b10110110010001010101000001111011;
		#400 //-9.686607e-20 * 3.294525e-14 = -2.9402133e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011101000111100011110111011100;
		b = 32'b00101111101101100001000011110100;
		correct = 32'b10101100110111101000000000101101;
		#400 //-2.0943106e-21 * 3.3117653e-10 = -6.32385e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110010011111110100010100111000;
		b = 32'b00001011010011011100001000101100;
		correct = 32'b11100110100111101100110100000000;
		#400 //-1.4858692e-08 * 3.9627643e-32 = -3.7495774e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111000010001000111001011000110;
		b = 32'b01010100010011001001111110011101;
		correct = 32'b11100011011101011100010110110010;
		#400 //-1.5937782e+34 * 3515404800000.0 = -4.5336977e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000100011100000000100011100101;
		b = 32'b10101100100000000010000001110011;
		correct = 32'b00010111011011111100110000011011;
		#400 //-2.8215949e-36 * -3.6415814e-12 = 7.748268e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000001001100110110000101100100;
		b = 32'b11100001110010001100101100001111;
		correct = 32'b10011110111001001011001100101111;
		#400 //11.211277 * -4.629976e+20 = -2.4214548e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011101011001010010101101100001;
		b = 32'b10011000111100111101100110110000;
		correct = 32'b01000011111100001001011001110000;
		#400 //-3.0330324e-21 * -6.3033836e-24 = 481.1753
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010000111111101010111100000111;
		b = 32'b00011110111000110100101001011101;
		correct = 32'b01110001100011110110110100111001;
		#400 //34183068000.0 * 2.4065316e-20 = 1.4204288e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001001001010001110010110101100;
		b = 32'b11100000111001110000001001000111;
		correct = 32'b00100111101110110010101100111010;
		#400 //-691802.75 * -1.3316756e+20 = 5.1949793e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010111001000111111100011000011;
		b = 32'b11001110001010101100001010101000;
		correct = 32'b11001000011101011101001010010111;
		#400 //180288820000000.0 * -716220900.0 = -251722.36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110010000100000110000010101101;
		b = 32'b11101100101011110001001001001011;
		correct = 32'b11000100110100110001111000011111;
		#400 //2.8596938e+30 * -1.6931872e+27 = -1688.9413
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101111010110110001110000011010;
		b = 32'b11011011010111111111111011101011;
		correct = 32'b11010011011110100110101001111000;
		#400 //6.781119e+28 * -6.3049205e+16 = -1075528100000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110101110111100100110100110011;
		b = 32'b11010011011000011100111111111100;
		correct = 32'b01100001111111000000010100010000;
		#400 //-5.636014e+32 * -969857040000.0 = 5.8111804e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111011000011100110111100001010;
		b = 32'b01010110011001001011111000011011;
		correct = 32'b01100100000111110110100000001011;
		#400 //7.395583e+35 * 62876287000000.0 = 1.1762118e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011111100111010110101101000011;
		b = 32'b00111010010110000100000011100010;
		correct = 32'b00100100101110100101101000011100;
		#400 //6.6669536e-20 * 0.00082494144 = 8.081729e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011000101001010001010000011110;
		b = 32'b10001111000111000000111101001000;
		correct = 32'b11001001000001110110010110110100;
		#400 //4.2671814e-24 * -7.694337e-30 = -554587.25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110100110001010010100001011101;
		b = 32'b10111101011100010100011000001100;
		correct = 32'b10110110110100010011000011111111;
		#400 //3.6723478e-07 * -0.058904693 = -6.2343893e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110010000010110101000110100011;
		b = 32'b10010110111110010101000110010111;
		correct = 32'b11011010100011110000110101101001;
		#400 //8.109427e-09 * -4.027961e-25 = -2.0132833e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001101101010011011000111000001;
		b = 32'b01001111101101011111010001100001;
		correct = 32'b10111101011011101100000000100001;
		#400 //-355874850.0 * 6105383400.0 = -0.058288697
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011010111000010011011100110;
		b = 32'b11001000111111000000011111101000;
		correct = 32'b01000001110111111001111001111000;
		#400 //-14427878.0 * -516159.25 = 27.952377
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100011101110101010100011111011;
		b = 32'b00011101010110001001100001010100;
		correct = 32'b01000101110111001001111001110111;
		#400 //2.0237726e-17 * 2.8666114e-21 = 7059.808
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111000011001010111001000110111;
		b = 32'b01101011010010100100000010011101;
		correct = 32'b10001100100100010011010111001111;
		#400 //-5.4704225e-05 * 2.4450814e+26 = -2.2373172e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101110011110010110111100011010;
		b = 32'b01111000100101001111011101010100;
		correct = 32'b10110101010101100101001111011101;
		#400 //-1.929902e+28 * 2.4171136e+34 = -7.984325e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000111001101110011100101110;
		b = 32'b00011011011010110001000100000100;
		correct = 32'b11010100111110110111011100111111;
		#400 //-1.6800408e-09 * 1.9444242e-22 = -8640299300000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100001111000110100001010101110;
		b = 32'b10111011011000101110001100111000;
		correct = 32'b01100110000000000011010111011011;
		#400 //-5.2402696e+20 * -0.0034620296 = 1.513641e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000111000100010100011101110111;
		b = 32'b10011001001100011101011111001011;
		correct = 32'b01101101010100010010000000010110;
		#400 //-37191.465 * -9.1942646e-24 = 4.0450723e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011101000010111001111110010011;
		b = 32'b10110011111100111100110011000001;
		correct = 32'b01101000100100101001110000111111;
		#400 //-6.288076e+17 * -1.1352814e-07 = 5.538782e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110100001100100000110010010000;
		b = 32'b10001111110010111000110001110000;
		correct = 32'b01100011110111111110110111111101;
		#400 //-1.6582112e-07 * -2.007144e-29 = 8.2615456e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111111000001111010000110011110;
		b = 32'b10111011100011111010110000111010;
		correct = 32'b01000010111100011010101111101010;
		#400 //-0.52980983 * -0.0043845447 = 120.83577
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011110100111010011100010011111;
		b = 32'b10111001010000000110011111110111;
		correct = 32'b00100100110100010010111110001111;
		#400 //-1.664644e-20 * -0.00018349277 = 9.071987e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111111000001010011101111100100;
		b = 32'b10111111000111101100101011110010;
		correct = 32'b11111111010101101100101110000101;
		#400 //1.770983e+38 * -0.6202842 = -2.8551152e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011110110001110110011011001101;
		b = 32'b01111111011101010001111111111101;
		correct = 32'b10011110110100000011111110000010;
		#400 //-7.1841985e+18 * 3.2582695e+38 = -2.2049123e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101101010100001001110011001100;
		b = 32'b01011010100110110110001000101000;
		correct = 32'b01010010001010111101100100110011;
		#400 //4.0351524e+27 * 2.1868273e+16 = 184520850000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001110011010101000110000010110;
		b = 32'b11100101001111011011000001111000;
		correct = 32'b10101000100111100100010100000001;
		#400 //983762300.0 * -5.598641e+22 = -1.757145e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010001010101110000111101001110;
		b = 32'b10110110000011101100101011101001;
		correct = 32'b11011010110000001100011111011000;
		#400 //57729670000.0 * -2.1277758e-06 = -2.7131463e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110100010101110011010110011100;
		b = 32'b01001101001011111000010001110000;
		correct = 32'b00100110100111001111001001000100;
		#400 //2.0042938e-07 * 184043260.0 = 1.0890341e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100110010100001101011101100110;
		b = 32'b10101000000011100010101000101100;
		correct = 32'b10111101101111000000100010000100;
		#400 //7.2456416e-16 * -7.891728e-15 = -0.09181312
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100110100000010100000000110;
		b = 32'b10010111011101100110011100110011;
		correct = 32'b11101100110110000100001101111011;
		#400 //1665.2507 * -7.9617143e-25 = -2.0915732e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101011110100100010000011111100;
		b = 32'b10010001000111101011101010111000;
		correct = 32'b01011010001010010111001011100001;
		#400 //-1.4930552e-12 * -1.252154e-28 = 1.1923895e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110110111111000000001010010000;
		b = 32'b10100000010010111011110000111000;
		correct = 32'b11010110000111100101010001010101;
		#400 //7.5104836e-06 * -1.7257045e-19 = -43521260000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001100111010101111010110101110;
		b = 32'b10100101001101100100101101111000;
		correct = 32'b10100111001001001111101010101001;
		#400 //3.6201272e-31 * -1.5811553e-16 = -2.2895455e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110000001000110110111011011011;
		b = 32'b01001110111101010101011111001010;
		correct = 32'b01100000101010101000100000111011;
		#400 //2.023203e+29 * 2058085600.0 = 9.830509e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110110100110101011000101001010;
		b = 32'b01111000000111011010011011100111;
		correct = 32'b00111101111110110011000111000100;
		#400 //1.5687687e+33 * 1.2790247e+34 = 0.122653514
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010011000100110000100001100001;
		b = 32'b01000011000000110111001001100101;
		correct = 32'b11001111100011110010110101011011;
		#400 //-631500770000.0 * 131.44685 = -4804228600.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101111101111011100000001011001;
		b = 32'b01000001110110000110000011110101;
		correct = 32'b01101101011000000111111100110010;
		#400 //1.174504e+29 * 27.047342 = 4.3424007e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011100011000110110000011110111;
		b = 32'b00110111010010011110001100101111;
		correct = 32'b10100100100100000010100101110100;
		#400 //-7.5233324e-22 * 1.2033429e-05 = -6.252027e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100110011110010111101100010111;
		b = 32'b00010111110010101100000110001010;
		correct = 32'b01001110000111010111111101010110;
		#400 //8.6556047e-16 * 1.31028e-24 = 660592000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101101011010000101111010110110;
		b = 32'b01001100111111110000000011110001;
		correct = 32'b01011111111010010100011100100010;
		#400 //4.4946888e+27 * 133695370.0 = 3.3618883e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110010110000110000100010010111;
		b = 32'b01011111001010100001100100000000;
		correct = 32'b10010011000100101100001110110101;
		#400 //-2.2704894e-08 * 1.2256828e+19 = -1.8524282e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000000000111001011100111011010;
		b = 32'b00001000010110101001011010110000;
		correct = 32'b01110111001101111000110010110010;
		#400 //2.4488435 * 6.577912e-34 = 3.722828e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011111110011100011111111111101;
		b = 32'b00011110101111001111111110111100;
		correct = 32'b11000000100010111010111011101011;
		#400 //-8.7350253e-20 * 2.0011044e-20 = -4.3651023
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111010101110101101100000110111;
		b = 32'b11011001000010100010011001100000;
		correct = 32'b10100001001011010001110111111001;
		#400 //0.0014255111 * -2430358800000000.0 = -5.865435e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001101101001001011111000011001;
		b = 32'b10000100011010111000001111000110;
		correct = 32'b01001000101100110001001001101111;
		#400 //-1.0153045e-30 * -2.7684625e-36 = 366739.47
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010011001110001101110011011110;
		b = 32'b00111001101101001101101101011011;
		correct = 32'b11011001000000101101010111001100;
		#400 //-793979500000.0 * 0.00034495708 = -2301676200000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101100110110111001011010000111;
		b = 32'b11100000010001011111010101000010;
		correct = 32'b00001100000011011111110001101000;
		#400 //-6.2410663e-12 * -5.705752e+19 = 1.0938201e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011011100101101100010001110011;
		b = 32'b01000101111000100011110000001001;
		correct = 32'b00010101001010101001101010001101;
		#400 //2.494237e-22 * 7239.5044 = 3.4453146e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011100001011001001101101001101;
		b = 32'b11011000110100101011100001010101;
		correct = 32'b10000010110100011011001001011100;
		#400 //5.711075e-22 * -1853513100000000.0 = -3.0812163e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011111001010010000100110110110;
		b = 32'b11010011101010001011111110100011;
		correct = 32'b00001011000000000011100000110000;
		#400 //-3.5795175e-20 * -1449539300000.0 = 2.4694174e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011100011000101011110111000;
		b = 32'b01110010111001101001011000000101;
		correct = 32'b10011000000110111100111101111100;
		#400 //-18394992.0 * 9.134453e+30 = -2.0138033e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101010010110100110000101011100;
		b = 32'b11001100001111000000011000010100;
		correct = 32'b11011101100101001010101001101011;
		#400 //6.60014e+25 * -49289296.0 = -1.3390615e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011111000010011000110111000011;
		b = 32'b01001110100100010101111011100101;
		correct = 32'b10001111111100100011101111111001;
		#400 //-2.912814e-20 * 1219457700.0 = -2.3886143e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100101010110011010010000110000;
		b = 32'b01110110000110111010111001110010;
		correct = 32'b10101110101100101111000101100101;
		#400 //-6.423639e+22 * 7.893986e+32 = -8.137383e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001010101001011010100100011011;
		b = 32'b01100010100000111101001110111010;
		correct = 32'b00100111101000001101100111101110;
		#400 //5428365.5 * 1.21589e+21 = 4.46452e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011100010101010001100110100110;
		b = 32'b01000001101111111101011000011110;
		correct = 32'b11011010000011100011000000011110;
		#400 //-2.3992948e+17 * 23.97955 = -1.0005588e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001010111000110001010100000111;
		b = 32'b10101100000001111010010110111110;
		correct = 32'b10011110010101100100011110100110;
		#400 //2.1867214e-32 * -1.927666e-12 = -1.1343882e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010101000110101010000001111010;
		b = 32'b10110011101000001001011100001001;
		correct = 32'b10100000111101100111111001111011;
		#400 //3.1226646e-26 * -7.478054e-08 = -4.175772e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001000111000101100000100010011;
		b = 32'b10011011111010110100111011010111;
		correct = 32'b00101100011101101011000110101101;
		#400 //-1.3647272e-33 * -3.8928438e-22 = 3.5057332e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010000000111100010010011110110;
		b = 32'b11111000000010001011010010011100;
		correct = 32'b00010111100101000001001011011001;
		#400 //-10612890000.0 * -1.1090868e+34 = 9.569034e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101100000011011100011101011000;
		b = 32'b11010011111111101000011011111111;
		correct = 32'b10010111100011101001100101011000;
		#400 //2.0147963e-12 * -2186373100000.0 = -9.215244e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111111011001000100111010011001;
		b = 32'b01011011101100011000111110101011;
		correct = 32'b11100011001001001001010011100001;
		#400 //-3.0347209e+38 * 9.995807e+16 = -3.035994e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111101100110100001100100010010;
		b = 32'b11101100011001111010000010011101;
		correct = 32'b11010000101010100101000000001000;
		#400 //2.560391e+37 * -1.12008136e+27 = -22858973000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000001111001010010101001001001;
		b = 32'b00001001110011001010000000110001;
		correct = 32'b00110111100011110101100110100111;
		#400 //8.418199e-38 * 4.9261857e-33 = 1.7088676e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001110000010001100000111011101;
		b = 32'b00101001010110010001011110110111;
		correct = 32'b10100100001000010100010001010110;
		#400 //-1.6856636e-30 * 4.820425e-14 = -3.4969193e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010000000110000011110101000100;
		b = 32'b10000011010011110100000100010011;
		correct = 32'b11001100001111000000101110110101;
		#400 //3.0023912e-29 * -6.0906534e-37 = -49295060.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110101111110100101111100011111;
		b = 32'b11100101001101000011011010110101;
		correct = 32'b01010000001100011101010010110100;
		#400 //-6.3476733e+32 * -5.3189696e+22 = 11934028000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011110100001000001010100100000;
		b = 32'b10111110110011010110110011100101;
		correct = 32'b00011111001001001001100110111100;
		#400 //-1.398478e-20 * -0.40122142 = 3.4855517e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010100100111101010101110100100;
		b = 32'b10001100010101100111101011101010;
		correct = 32'b01000111101111010110001011110001;
		#400 //-1.6021623e-26 * -1.6522948e-31 = 96965.88
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101000101010100000101000001011;
		b = 32'b00111000000001101010010101000100;
		correct = 32'b00110000001000011010010110010011;
		#400 //1.8878147e-14 * 3.2102005e-05 = 5.8806754e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001000110000110000000101000001;
		b = 32'b01011111010101110110110100110011;
		correct = 32'b10101000111001111011101101101100;
		#400 //-399370.03 * 1.552312e+19 = -2.5727433e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000000011101010000001100100101;
		b = 32'b01110000001110011100101110110101;
		correct = 32'b10001111101010001100101111000101;
		#400 //-3.828317 * 2.3000397e+29 = -1.6644568e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111100111000000110111110010101;
		b = 32'b00000001111100011100001011001011;
		correct = 32'b11111010011011011010011110010001;
		#400 //-0.027396956 * 8.880893e-38 = -3.0849325e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110011010001001000111110100000;
		b = 32'b11010011110000001111000100100000;
		correct = 32'b11011111000000100110011010100111;
		#400 //1.557317e+31 * -1657358300000.0 = -9.396381e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001001110000100100101010101110;
		b = 32'b10110010010111000110001100010010;
		correct = 32'b11010110111000011011000000011011;
		#400 //1591637.8 * -1.2828211e-08 = -124073240000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100100010000100001100111011111;
		b = 32'b01001011100001010011111010100110;
		correct = 32'b00011000001110100111011000000000;
		#400 //4.2088958e-17 * 17464652.0 = 2.4099511e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001100110100011100000000110011;
		b = 32'b10000011100011111110111101011011;
		correct = 32'b01001000101110101000011110000100;
		#400 //-3.2317224e-31 * -8.459738e-37 = 382012.12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100011000001000101111111110000;
		b = 32'b10101011100101000001010110101001;
		correct = 32'b11110110111001001101011101111011;
		#400 //2.4418832e+21 * -1.0522044e-12 = -2.3207308e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010110100111010111001000110000;
		b = 32'b01111110100111001011001011010100;
		correct = 32'b10010111100000001001110001010000;
		#400 //-86556880000000.0 * 1.0414405e+38 = -8.311265e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011001011110000011000001001010;
		b = 32'b00111000010101100101000000100001;
		correct = 32'b01100000100101000011101110000011;
		#400 //4366180500000000.0 * 5.10962e-05 = 8.54502e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000001011001010100101000100001;
		b = 32'b00001101111101101101110011111110;
		correct = 32'b10110010111011011100011010100001;
		#400 //-4.2113842e-38 * 1.5214122e-30 = -2.7680757e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001101011011001111100111011011;
		b = 32'b00100010000001010001110110100111;
		correct = 32'b10101010111000111101111001100010;
		#400 //-7.3023867e-31 * 1.8040559e-18 = -4.047761e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100011000000110011000111011010;
		b = 32'b00111000100110000100001101001001;
		correct = 32'b11101001110111001001010000000001;
		#400 //-2.4201157e+21 * 7.260458e-05 = -3.3332826e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011000010001101000100101111010;
		b = 32'b00011000111100110111000001001101;
		correct = 32'b00111110110100001100100000001100;
		#400 //2.5660308e-24 * 6.2927423e-24 = 0.40777624
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111001001111101101011011101001;
		b = 32'b01010111000111110010110011010010;
		correct = 32'b10100001100110010111011001111011;
		#400 //-0.00018199872 * 175014850000000.0 = -1.0399045e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100100111100010011010010010011;
		b = 32'b01011101101011100011110010111011;
		correct = 32'b01000110101100010011001001100100;
		#400 //3.559563e+22 * 1.5693894e+18 = 22681.195
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000001000101111010110011001010;
		b = 32'b01000000000000001011000000010111;
		correct = 32'b10000000100101101101110100111111;
		#400 //-2.785829e-38 * 2.0107477 = -1.3854693e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001101110000110001010101000111;
		b = 32'b00111011010010101100100001110110;
		correct = 32'b10010001111101100100011110000011;
		#400 //-1.2022925e-30 * 0.0030942238 = -3.885603e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000011101000111010010000110100;
		b = 32'b11100101001101101011000101111001;
		correct = 32'b00011101111001010100110110110010;
		#400 //-327.28284 * -5.392153e+22 = 6.069613e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010000101010011111111000010;
		b = 32'b11101100111011110001110110110000;
		correct = 32'b00001100100111111100100110011110;
		#400 //-0.00056933996 * -2.3125877e+27 = 2.4619173e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101110110000110100010011001011;
		b = 32'b01000111100111011011010101110011;
		correct = 32'b10100110100111100111110000001000;
		#400 //-8.8797934e-11 * 80746.9 = -1.0997071e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101000010011110110100010111010;
		b = 32'b11001110011000111000011001011100;
		correct = 32'b10011001011010010101110111100010;
		#400 //1.1513517e-14 * -954308350.0 = -1.2064777e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011000010111000110000011011110;
		b = 32'b10000000101010010111101011000010;
		correct = 32'b11010111001001100111000100001001;
		#400 //2.8483239e-24 * -1.5564236e-38 = -183004410000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000000100110010110100001000110;
		b = 32'b01011101010100001101111111001100;
		correct = 32'b10100010101111000000010011001111;
		#400 //-4.7939787 * 9.406858e+17 = -5.0962593e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011010100000010111000100001111;
		b = 32'b01010101000000011111100100101010;
		correct = 32'b10000100111111101111001111101100;
		#400 //-5.3535806e-23 * 8931697000000.0 = -5.993912e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010101001110001110001100011101;
		b = 32'b10100011011011101100110001001011;
		correct = 32'b11110001010001100011010010100101;
		#400 //12705349000000.0 * -1.29452666e-17 = -9.814668e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011011000001111110010010011;
		b = 32'b11011001000110011110010001101000;
		correct = 32'b00110001101110110010001000000010;
		#400 //-14744723.0 * -2707300400000000.0 = 5.4462825e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100110000100110110010101010111;
		b = 32'b10001000010110011111100011000011;
		correct = 32'b01011101001011010001110001110101;
		#400 //-5.113821e-16 * -6.559348e-34 = 7.7962336e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010011111001100111100000111110;
		b = 32'b00111101101100110010000111111100;
		correct = 32'b11010101101001001010111011011010;
		#400 //-1979719600000.0 * 0.087467164 = -22633861000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011111000110011001100100110011;
		b = 32'b01011000010111011010110111100110;
		correct = 32'b11000110001100010110000011110111;
		#400 //-1.1067934e+19 * 974955800000000.0 = -11352.241
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111101110000011000010011110101;
		b = 32'b01000111101111101101101001010110;
		correct = 32'b00110101100000011100100111010001;
		#400 //0.09449188 * 97716.67 = 9.669985e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111010111111111011000101010110;
		b = 32'b01100011011110111111100010101001;
		correct = 32'b00010111000000011110001111110100;
		#400 //0.0019507806 * 4.6480506e+21 = 4.1969865e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000000111100110110010100111110;
		b = 32'b10101110100000101101111110000010;
		correct = 32'b01010001111011100000110101011100;
		#400 //-7.6061087 * -5.9514185e-11 = 127803290000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111011111101001111101111100111;
		b = 32'b00011101101011110010011010010101;
		correct = 32'b01011101101100110000100010111011;
		#400 //0.007476318 * 4.6362007e-21 = 1.6125958e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001010011011011100111101111100;
		b = 32'b10010010011110100011000111101101;
		correct = 32'b01110111011100110101010000000000;
		#400 //-3896287.0 * -7.894763e-28 = 4.9352807e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110111101011100011010110001100;
		b = 32'b01110000011000110100001100111011;
		correct = 32'b01000110110001000011110011101001;
		#400 //7.0667634e+33 * 2.813375e+29 = 25118.455
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100101111001000000011000001;
		b = 32'b10101001011011010011101100000101;
		correct = 32'b11011010110010110110101011001000;
		#400 //1508.0236 * -5.2675763e-14 = -2.8628414e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010010010000110100010100111100;
		b = 32'b00000011110111101011110011001010;
		correct = 32'b01001101111000000110111001100011;
		#400 //6.161649e-28 * 1.3091331e-36 = 470666340.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111111110011101011011101000000;
		b = 32'b01011010110100001100101110100101;
		correct = 32'b10100100011111010111001100111110;
		#400 //-1.6149673 * 2.9385352e+16 = -5.4958244e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101010101010001011010111000011;
		b = 32'b11100100100000110100111000000100;
		correct = 32'b11000101101001000111011010111101;
		#400 //1.0197894e+26 * -1.937716e+22 = -5262.8423
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001110110010000110111110001110;
		b = 32'b10101110100101110100111000000011;
		correct = 32'b11011111101010011001000001001001;
		#400 //1681377000.0 * -6.880543e-11 = -2.4436692e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110010000010110100110101101000;
		b = 32'b11000000000100110110001100010101;
		correct = 32'b01110001011100011111010100100010;
		#400 //-2.7591677e+30 * -2.3029225 = 1.19811576e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010011100011001001011011011100;
		b = 32'b01000011100100101000010000100010;
		correct = 32'b11001111011101011010010011110011;
		#400 //-1207652800000.0 * 293.0323 = -4121228000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101001101000000111110001000011;
		b = 32'b11011100101001010101100011011010;
		correct = 32'b10001100011110000111100100001110;
		#400 //7.126983e-14 * -3.723285e+17 = -1.9141654e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011100000001110001001011111000;
		b = 32'b00110010101000000111001010010100;
		correct = 32'b00101000110101111000010000000100;
		#400 //4.469227e-22 * 1.8678556e-08 = 2.3927048e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111000111000110101000001100010;
		b = 32'b11100000110111101111101001110001;
		correct = 32'b10010111100000100111110100101001;
		#400 //0.00010839176 * -1.2853823e+20 = -8.432648e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101101111000111100100111011111;
		b = 32'b11101110011000011110111011011001;
		correct = 32'b00111111000000010000110100011111;
		#400 //-8.812143e+27 * -1.7480719e+28 = 0.50410646
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011100000100010110010110000000;
		b = 32'b01111001110100000000010111010101;
		correct = 32'b00100001101100101110111000001111;
		#400 //1.6370189e+17 * 1.350145e+35 = 1.2124763e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101011010101100010000100110000;
		b = 32'b00010111110011011011101111111000;
		correct = 32'b01010011000001010011100100101001;
		#400 //7.607413e-13 * 1.3295264e-24 = 572189640000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011001111001110111001111010010;
		b = 32'b10100010000111001001101100000010;
		correct = 32'b01110111001111010010110011101000;
		#400 //-8143508000000000.0 * -2.1224003e-18 = 3.8369333e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100001011100000110011110100010;
		b = 32'b10100111101000100011100010010101;
		correct = 32'b01111001001111011011000011010000;
		#400 //-2.7716788e+20 * -4.502538e-15 = 6.1558143e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100011100000111100001001011111;
		b = 32'b10101111011100011100100111101010;
		correct = 32'b01110011100010111000000011100101;
		#400 //-4.861059e+21 * -2.1990557e-10 = 2.210521e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101001110011101010001000111001;
		b = 32'b11110111010011010101111111011000;
		correct = 32'b10110010000000001100100011101100;
		#400 //3.12256e+25 * -4.1654875e+33 = -7.496265e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001001011110001101101000001110;
		b = 32'b10001100000000101111101001001101;
		correct = 32'b01111100111100110011000110111000;
		#400 //-1019296.9 * -1.0090158e-31 = 1.01018924e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101101110000100001001100110011;
		b = 32'b11011100101110101010011000111100;
		correct = 32'b10010000100001010001011110100100;
		#400 //2.2063773e-11 * -4.2029698e+17 = -5.2495674e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100010110111111100111000000000;
		b = 32'b01111111010010111101101001011001;
		correct = 32'b10100011000011001000011100011101;
		#400 //-2.0642339e+21 * 2.70967e+38 = -7.6180266e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000111000001001000010000101011;
		b = 32'b00111001000000000010000101101010;
		correct = 32'b00001101100001000110000110011100;
		#400 //9.969417e-35 * 0.00012219479 = 8.158627e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101011101101000110001010010001;
		b = 32'b00001110001111001001000110010111;
		correct = 32'b11011100111101001110001111001110;
		#400 //-1.2817127e-12 * 2.3242888e-30 = -5.5144295e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110010010111001011111010111111;
		b = 32'b01100010100110011111101111000101;
		correct = 32'b01001111001101110111111100000011;
		#400 //4.3723072e+30 * 1.4202469e+21 = 3078554400.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101000100011110101111101100000;
		b = 32'b01010100001000101110101111010110;
		correct = 32'b00010011111000010100100001101111;
		#400 //1.5917552e-14 * 2798965500000.0 = 5.686941e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111011100111000001000101100111;
		b = 32'b00111111001000101100000011101011;
		correct = 32'b00111011111101010111101111101000;
		#400 //0.0047628167 * 0.6357562 = 0.0074915774
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011101011001011011000010010010;
		b = 32'b00010011110000000000100001001011;
		correct = 32'b11001001000110010001100111000100;
		#400 //-3.0399182e-21 * 4.847579e-27 = -627100.25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011011010101000101111010000100;
		b = 32'b00011110010101001001000000001100;
		correct = 32'b01111100011111111100010001011001;
		#400 //5.9776616e+16 * 1.1252975e-20 = 5.3120724e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101010010101100111000101000011;
		b = 32'b00110011010100010010101010011011;
		correct = 32'b10110110100000110011101010001010;
		#400 //-1.9046314e-13 * 4.8700354e-08 = -3.910919e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010011100110000011100110001010;
		b = 32'b01011000011000011001001111000000;
		correct = 32'b10111010101011001100000100111100;
		#400 //-1307600700000.0 * 992098800000000.0 = -0.0013180147
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111110110010101001010000011011;
		b = 32'b01111101000101101100100110001101;
		correct = 32'b11000001001010111111011011100101;
		#400 //-1.3463653e+38 * 1.252692e+37 = -10.747777
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011110000110110010000110100000;
		b = 32'b00100001001110010011010110111001;
		correct = 32'b00111100010101100110110011001110;
		#400 //8.212585e-21 * 6.275154e-19 = 0.0130874645
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000000110101101001010101010010;
		b = 32'b00111011000000000010101011111011;
		correct = 32'b10000101010101100100110101011100;
		#400 //-1.9706362e-38 * 0.0019556868 = -1.007644e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000111111010111011001010111110;
		b = 32'b00100111101011000001010001000110;
		correct = 32'b10011111101011110101001010010110;
		#400 //-3.5463925e-34 * 4.776157e-15 = -7.425201e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100101101001011111101101010101;
		b = 32'b10101101100111101110011011110100;
		correct = 32'b00110111100001011011001111101100;
		#400 //-2.8793247e-16 * -1.8065084e-11 = 1.5938618e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101110100011111001011011101000;
		b = 32'b00110011011110111111111010000010;
		correct = 32'b01111010100100011101111100111111;
		#400 //2.2219395e+28 * 5.8671965e-08 = 3.787055e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100011001100100100110011111001;
		b = 32'b01010000101101101111010011000111;
		correct = 32'b00010001111110010111110001100000;
		#400 //9.665699e-18 * 24555960000.0 = 3.9361925e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101011010011000100110000001110;
		b = 32'b11010010101111000111000011000001;
		correct = 32'b11011000000010101100010101010010;
		#400 //2.4698003e+26 * -404672770000.0 = -610320360000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010001110101111011110000110110;
		b = 32'b11111000100001010011010110110000;
		correct = 32'b10011000110011110100110001001001;
		#400 //115821950000.0 * -2.1614512e+34 = -5.3585274e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100010111001101100111101000000;
		b = 32'b00111110111011101000000101100001;
		correct = 32'b01100011011101111011110101011100;
		#400 //2.1288425e+21 * 0.46583083 = 4.5699906e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111101010110110010100010000111;
		b = 32'b00110010011101100011101001011111;
		correct = 32'b11001010011000111101101100100010;
		#400 //-0.053505447 * 1.4332357e-08 = -3733192.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000110101110111000001101000011;
		b = 32'b11110101111000111110110110101111;
		correct = 32'b00010000010100101001101101010001;
		#400 //-24001.63 * -5.7786728e+32 = 4.153485e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111110111100100010001011101000;
		b = 32'b11111100100000010000110110010100;
		correct = 32'b11000001111100000010100100011100;
		#400 //1.6092721e+38 * -5.3606535e+36 = -30.020073
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010001011000011011001001101110;
		b = 32'b00111101010000001000011100101000;
		correct = 32'b00010011100101100000110101010011;
		#400 //1.7804353e-28 * 0.047003895 = 3.7878462e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000101011110011100000000100010;
		b = 32'b00111000001001101000011001010000;
		correct = 32'b00001100101111111111100011010011;
		#400 //1.1743213e-35 * 3.9702572e-05 = 2.9577965e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110001001111111000100100000101;
		b = 32'b01001011001001100010100011111010;
		correct = 32'b11100101100100111000110000101100;
		#400 //-9.484365e+29 * 10889466.0 = -8.70967e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001100110100010100100101010101;
		b = 32'b10011010010111110000001101010001;
		correct = 32'b11110001111100000011111000111110;
		#400 //109726376.0 * -4.6117998e-23 = -2.3792528e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010110000110110010001100001111;
		b = 32'b10011010001110111010110101011110;
		correct = 32'b01111011010100111001110100010111;
		#400 //-42643720000000.0 * -3.881074e-23 = 1.0987608e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100010010101001011111001110110;
		b = 32'b01001001001011111110111100001111;
		correct = 32'b00011000100110101100011111110110;
		#400 //2.8832187e-18 * 720624.94 = 4.0009976e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101010001101110010000011000000;
		b = 32'b10101000010101001110110000001001;
		correct = 32'b11000001010111000010110110010100;
		#400 //1.6265028e-13 * -1.1819546e-14 = -13.761127
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011011010001001100101010011110;
		b = 32'b10011101000101010000111100110110;
		correct = 32'b01111101101010001111110100000110;
		#400 //-5.5391875e+16 * -1.972785e-21 = 2.807801e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000011000101110111000111010;
		b = 32'b01011011000000110100111010010110;
		correct = 32'b10010100110111010011011100011110;
		#400 //-8.255686e-10 * 3.695963e+16 = -2.2337037e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110101001000100100000010011000;
		b = 32'b01111101010100100000010101010100;
		correct = 32'b10110111010001011100011000010001;
		#400 //-2.0567925e+32 * 1.7447847e+37 = -1.1788231e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011001000000111011010100110;
		b = 32'b01111110011011010110011011000111;
		correct = 32'b10001100001011010000100011010110;
		#400 //-10516134.0 * 7.889017e+37 = -1.3330094e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100011001101101010010000101101;
		b = 32'b01000110010101010101011000001011;
		correct = 32'b10011100010110110010101010101111;
		#400 //-9.901005e-18 * 13653.511 = -7.251619e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110110011011100011000011011010;
		b = 32'b01000010101000100000100001000000;
		correct = 32'b00110011001111000010100110101001;
		#400 //3.54932e-06 * 81.01611 = 4.381005e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001010011001100111110110010011;
		b = 32'b01011111001010010000111111101100;
		correct = 32'b10101010101011101000001000101100;
		#400 //-3776356.8 * 1.2182215e+19 = -3.0998934e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101101101100011100011001101110;
		b = 32'b11010100011000011100011000111110;
		correct = 32'b00011000110010011001001100100111;
		#400 //-2.021069e-11 * -3878774400000.0 = 5.210587e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101111100101000111001011011101;
		b = 32'b00001111110000100110011110000100;
		correct = 32'b01011111010000110111101111001101;
		#400 //2.7002658e-10 * 1.916975e-29 = 1.4086078e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101110111110100101100100010001;
		b = 32'b10110010011111010110111111010111;
		correct = 32'b00111011111111001110000100111011;
		#400 //-1.1384505e-10 * -1.4751968e-08 = 0.0077172793
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100110001110101101010111011110;
		b = 32'b10101110111011010101001001110110;
		correct = 32'b11110110110010011000101000110101;
		#400 //2.2057633e+23 * -1.079216e-10 = -2.0438571e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101000100010101010011101101100;
		b = 32'b11101101111111001001101111110100;
		correct = 32'b10111010000011001000001111100010;
		#400 //5.2381997e+24 * -9.772345e+27 = -0.0005360228
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000010011010010111000000011001;
		b = 32'b01010000010110110101110111000110;
		correct = 32'b00110001100010000011010111110100;
		#400 //58.35947 * 14721423000.0 = 3.9642547e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010111000110111111000111110101;
		b = 32'b10010101010010001011111001011101;
		correct = 32'b11000001010001101101111011010001;
		#400 //5.0388594e-25 * -4.053985e-26 = -12.429399
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001010111011001100010101111100;
		b = 32'b01100001110001001000011111010010;
		correct = 32'b10101000100110100011010101110101;
		#400 //-7758526.0 * 4.531686e+20 = -1.7120618e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001001011001100001110100111001;
		b = 32'b10110110011011110111111101110110;
		correct = 32'b01010010011101011111100000111110;
		#400 //-942547.56 * -3.5687967e-06 = 264107950000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110011010001110000011010111000;
		b = 32'b10000100011100001010000001000000;
		correct = 32'b11101110010100111011111000001101;
		#400 //4.633941e-08 * -2.8285448e-36 = -1.6382774e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010111101000111100100000011110;
		b = 32'b01001111000000111110110010110101;
		correct = 32'b10001000000111101110100011001011;
		#400 //-1.0584145e-24 * 2213328100.0 = -4.7820042e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001010010100111001010100000100;
		b = 32'b10110001110100111011100001000000;
		correct = 32'b10010111111111111101010101100110;
		#400 //1.0187307e-32 * -6.161855e-09 = -1.6532858e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011001001000110011001001000001;
		b = 32'b11000010010111111110001101000101;
		correct = 32'b11010110001110101001101010000011;
		#400 //2870979700000000.0 * -55.971943 = -51293196000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001110111100011010010111110011;
		b = 32'b01101000001011001000001001101010;
		correct = 32'b10100110001100110100110011011010;
		#400 //-2027092400.0 * 3.258611e+24 = -6.2207254e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000010110110110001110100000100;
		b = 32'b10101000001001000010110000011111;
		correct = 32'b00011010001010101101010111110100;
		#400 //-3.2195812e-37 * -9.113396e-15 = 3.5328006e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110100100111110011010111010001;
		b = 32'b10000111001110001001010100010001;
		correct = 32'b11101100110111001100111110100011;
		#400 //2.9655214e-07 * -1.3886428e-34 = -2.1355537e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110010100100110100111100111000;
		b = 32'b01101000110011111100001011111001;
		correct = 32'b10001001001101011000001100010000;
		#400 //-1.7149077e-08 * 7.849012e+24 = -2.1848708e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010111000101001000101011100101;
		b = 32'b01110100000011100111000000010001;
		correct = 32'b10100010100001010111110001101011;
		#400 //-163324270000000.0 * 4.514033e+31 = -3.6181455e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101100111111011010101010010011;
		b = 32'b00110000000011011101101100011101;
		correct = 32'b00111100011001001110001110100011;
		#400 //7.20963e-12 * 5.160688e-10 = 0.013970288
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100100101001110111110001000011;
		b = 32'b11011010100100010101100010001101;
		correct = 32'b10001001100100110111111101010000;
		#400 //7.263521e-17 * -2.0455617e+16 = -3.5508687e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101000011100010101000010011100;
		b = 32'b01000001110100100011100011011010;
		correct = 32'b10100110000100101110111010001001;
		#400 //-1.3395667e-14 * 26.27776 = -5.09772e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011011000101001010010011010010;
		b = 32'b11101110101101100000110000111000;
		correct = 32'b00101011110100010000011011010000;
		#400 //-4.183952e+16 * -2.8170522e+28 = 1.4852234e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110010110000001000011101110100;
		b = 32'b11100000010010101000100000101101;
		correct = 32'b00010001111100110101101101000000;
		#400 //-2.2413339e-08 * -5.8375856e+19 = 3.8394877e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001101110100101001101010110110;
		b = 32'b00000011100100001011010001010000;
		correct = 32'b01001001101110100100101011101011;
		#400 //1.29794945e-30 * 8.504957e-37 = 1526109.4
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010100011000101110000100000110;
		b = 32'b11010011001111000111010100001100;
		correct = 32'b11000000100110100001100010010111;
		#400 //3897751500000.0 * -809417600000.0 = -4.8155017
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010101101001000110001010000010;
		b = 32'b00111000011010111101011110100000;
		correct = 32'b10011100101100100110111101011001;
		#400 //-6.639449e-26 * 5.6229183e-05 = -1.1807835e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001000100001111101000010100111;
		b = 32'b00000110111111010101101001101110;
		correct = 32'b01000001000010010011101111100001;
		#400 //8.174071e-34 * 9.5300897e-35 = 8.577119
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100110100101101000001100100110;
		b = 32'b11001010000101111101101001010010;
		correct = 32'b00011011111111011011110101110111;
		#400 //-1.0443889e-15 * -2487956.5 = 4.1977778e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100110011001111000010100100;
		b = 32'b00100011111001100011110101111010;
		correct = 32'b01100000011000111101111010000101;
		#400 //1639.52 * 2.4962686e-17 = 6.567883e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010011011101110110000011100000;
		b = 32'b10101001111000110000111111011000;
		correct = 32'b11101001000010110111001111110001;
		#400 //1062482200000.0 * -1.00835735e-13 = -1.0536763e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010000110101101010001100011000;
		b = 32'b00011111111000000011101111111010;
		correct = 32'b01110000011101010000101100010001;
		#400 //28808102000.0 * 9.496691e-20 = 3.0334882e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100111000011010110011011000001;
		b = 32'b10111011111010100100110001111000;
		correct = 32'b11101010100110100111111110010001;
		#400 //6.6774915e+23 * -0.007150229 = -9.33885e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001111001101100110000010001101;
		b = 32'b10000111110110000010010000000000;
		correct = 32'b11000110110110000000001010010100;
		#400 //8.991888e-30 * -3.2521227e-34 = -27649.29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010101010101000000110100010100;
		b = 32'b00001111000111101110011010010011;
		correct = 32'b01000101101010101101000010000011;
		#400 //4.2823376e-26 * 7.8344084e-30 = 5466.064
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110011100100011110110101101000;
		b = 32'b11111101011001000010010011001010;
		correct = 32'b10110101101000111011111010111101;
		#400 //2.3123114e+31 * -1.8953438e+37 = -1.2199959e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110000111100110011100111010011;
		b = 32'b00111111110010000000101001101011;
		correct = 32'b01110000100110111010001000000101;
		#400 //6.021981e+29 * 1.5628179 = 3.8532837e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000101000000000101110011001101;
		b = 32'b10111111000001001100010111111111;
		correct = 32'b00000101011101110111111011001101;
		#400 //-6.035576e-36 * -0.5186462 = 1.1637174e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011000010110001001011011100110;
		b = 32'b10101110110001001010110001100101;
		correct = 32'b00101001000011001111011000111100;
		#400 //-2.799353e-24 * -8.9436715e-11 = 3.129982e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101000101110001001110001110000;
		b = 32'b11000100010011101000111000010001;
		correct = 32'b00100011111001001100110110100000;
		#400 //-2.0495948e-14 * -826.2198 = 2.4806895e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011110001111111110000100111100;
		b = 32'b11011110110100110001011011101010;
		correct = 32'b10111110111010001011010000001110;
		#400 //3.4565996e+18 * -7.605301e+18 = -0.4544987
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001010101101001100001110011011;
		b = 32'b00111010000100101100000001110111;
		correct = 32'b10010000000111011010101010001101;
		#400 //-1.7406948e-32 * 0.00055981375 = -3.1094178e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011110111011011010111000001101;
		b = 32'b10110100101101000101001010001110;
		correct = 32'b01101001101010001011011011101101;
		#400 //-8.5633204e+18 * -3.358768e-07 = 2.5495423e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000110110100010001110010010100;
		b = 32'b01001110010100011111101001001001;
		correct = 32'b10110111111111101111000110110011;
		#400 //-26766.29 * 880710200.0 = -3.039171e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010110110000010011000111000001;
		b = 32'b00000001101001001111011100111110;
		correct = 32'b11010100100101011110011100101111;
		#400 //-3.121223e-25 * 6.059886e-38 = -5150630000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011101110010110010100111000011;
		b = 32'b10001001100110011111001001000110;
		correct = 32'b11010011101010001110101111110011;
		#400 //5.3776833e-21 * -3.7061243e-33 = -1451026200000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011110010010100110011010101010;
		b = 32'b01001000100101111000000010111010;
		correct = 32'b01010101001010110000000010010110;
		#400 //3.6461328e+18 * 310277.8 = 11751188000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100111010001011100011100000100;
		b = 32'b11010011111011111110100100110101;
		correct = 32'b00010010110100110000101001110110;
		#400 //-2.7447129e-15 * -2060819500000.0 = 1.3318551e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011101010001101101101100111011;
		b = 32'b11100000111100100010000000100011;
		correct = 32'b00111011110100100100000001011011;
		#400 //-8.955695e+17 * -1.3957587e+20 = 0.006416363
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111111111101101000000100100010;
		b = 32'b00010110011000010010111011111101;
		correct = 32'b11101001000011000001111010001100;
		#400 //-1.9258158 * 1.8190182e-25 = -1.0587117e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110001010010101110110010111100;
		b = 32'b10001000101101001111001111000101;
		correct = 32'b11101000000011111000101011101101;
		#400 //2.9529437e-09 * -1.0890666e-33 = -2.7114445e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001110111111011011111100101101;
		b = 32'b10001110100011100101001011001101;
		correct = 32'b10111111111001000011010110101110;
		#400 //6.255341e-30 * -3.5085437e-30 = -1.7828882
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110010011010110000101100000100;
		b = 32'b11011001010101110011010001010111;
		correct = 32'b10011000100010111100110010110110;
		#400 //1.3681305e-08 * -3785916800000000.0 = -3.6137363e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101000110011100101101010000000;
		b = 32'b01011001011011010001101111111100;
		correct = 32'b10001110110111101100101100111011;
		#400 //-2.2909842e-14 * 4171271200000000.0 = -5.492293e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001110001100000000111100000000;
		b = 32'b01001011010001100111011111010001;
		correct = 32'b11000010011000110001100000110010;
		#400 //-738443260.0 * 13006801.0 = -56.77363
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000101010010000011111110100101;
		b = 32'b00100001111000110111110010001010;
		correct = 32'b10100010111000010101100100011101;
		#400 //-9.4156445e-36 * 1.5415084e-18 = -6.1080725e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001100100001010011000000000000;
		b = 32'b10010000000100011110010000110101;
		correct = 32'b10111011111010011011010101000010;
		#400 //2.0520784e-31 * -2.8772012e-29 = -0.0071322033
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110101111011101100011001000110;
		b = 32'b10000010010100110010111001101100;
		correct = 32'b11110011000100001011100110000000;
		#400 //1.7790087e-06 * -1.5515154e-37 = -1.1466265e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011111110110111000001110101001;
		b = 32'b11001111010000110100001110001000;
		correct = 32'b00010000000011111110010110010011;
		#400 //-9.296792e-20 * -3275982800.0 = 2.8378635e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010010000101111111111000101111;
		b = 32'b10011001000011000101110100101100;
		correct = 32'b00111000100010101001101011001000;
		#400 //-4.7960504e-28 * -7.256646e-24 = 6.609183e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101001101010001001101111101001;
		b = 32'b10010010010101111000011010100110;
		correct = 32'b11010110110010000100010110111110;
		#400 //7.487745e-14 * -6.8008005e-28 = -110100930000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000000111101011101000001111010;
		b = 32'b10001000110111100111101011100000;
		correct = 32'b01110111100011010110110011001111;
		#400 //-7.681699 * -1.3390027e-33 = 5.736881e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101001010001000000010100111110;
		b = 32'b01111111111011011100000001001010;
		correct = 32'b01111111111011011100000001001010;
		#400 //4.352529e-14 * nan = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100110000000101010011100101001;
		b = 32'b10110101010111001011011111111110;
		correct = 32'b00110000000101111000100110011001;
		#400 //-4.5329355e-16 * -8.222413e-07 = 5.512902e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111000110101000110110100001000;
		b = 32'b10100111110100101100110011010101;
		correct = 32'b01010000100000001111110010111000;
		#400 //-0.000101292564 * -5.850879e-15 = 17312367000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100000110100011000110011110111;
		b = 32'b00101001111010111010010001111000;
		correct = 32'b11110110011000111010011101110001;
		#400 //-1.2079772e+20 * 1.0464627e-13 = -1.1543433e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000101000000010100111100011011;
		b = 32'b01110110111100010110100001101011;
		correct = 32'b10001101100010010010000000001101;
		#400 //-2068.944 * 2.4481668e+33 = -8.450993e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010110010101110111010111111101;
		b = 32'b10100001101100110111100011011001;
		correct = 32'b00110100000110011010101011010111;
		#400 //-1.7404792e-25 * -1.21615e-18 = 1.4311387e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100000110111100011111010100010;
		b = 32'b11000110000100100001000111110111;
		correct = 32'b01011010010000101100000001000011;
		#400 //-1.2811532e+20 * -9348.491 = 1.3704385e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010000110010011011000101011000;
		b = 32'b00100110110010101001001001101110;
		correct = 32'b10101001011111101110001110001100;
		#400 //-7.955376e-29 * 1.4056256e-15 = -5.6596695e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010001011110011010010001111100;
		b = 32'b11001101001110001001010101000100;
		correct = 32'b11000011101011010001110110100100;
		#400 //67012903000.0 * -193549380.0 = -346.23157
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011010110111001010011111100011;
		b = 32'b10110111101000110101100101001111;
		correct = 32'b01100010101011001110011111011010;
		#400 //-3.1054544e+16 * -1.9472702e-05 = 1.5947733e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100110011011011100110000111101;
		b = 32'b00111110110010100010100001001000;
		correct = 32'b01100111000101101001000100000100;
		#400 //2.807421e+23 * 0.39483857 = 7.1103004e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001100100111000110111011110100;
		b = 32'b10100001101100010000000111011101;
		correct = 32'b10101010011000100011111010100011;
		#400 //2.4102383e-31 * -1.199448e-18 = -2.0094564e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011111000111001110000010111001;
		b = 32'b00011011101011110101110100110100;
		correct = 32'b11000010111001010000001101101110;
		#400 //-3.322017e-20 * 2.9011553e-22 = -114.5067
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001010001001100010011001011011;
		b = 32'b00110010001000111010000001001101;
		correct = 32'b10010111100000011111100101100100;
		#400 //-7.999823e-33 * 9.524297e-09 = -8.399385e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100100101111010111110001000011;
		b = 32'b10101010100011100011010100111010;
		correct = 32'b01111001101010101000110111010100;
		#400 //-2.796311e+22 * -2.52612e-13 = 1.1069589e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000111111100000011100101101000;
		b = 32'b10101000110100000001111111101110;
		correct = 32'b10011110100100111011110111100001;
		#400 //3.6144927e-34 * -2.3106486e-14 = -1.5642762e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101100010100010100010011101000;
		b = 32'b10000000110110001100010001001100;
		correct = 32'b01101010111101110010010100110111;
		#400 //-2.9738937e-12 * -1.9906885e-38 = 1.4939021e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100010100001111110101010010101;
		b = 32'b10010110110111011111100001100100;
		correct = 32'b01001011000111001100000011011011;
		#400 //-3.6840197e-18 * -3.5861232e-25 = 10272987.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000110100101000011010010100100;
		b = 32'b10000110110100010110011100110011;
		correct = 32'b00111111001101010010111101001000;
		#400 //-5.574876e-35 * -7.87687e-35 = 0.7077527
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010010110011011110010010110111;
		b = 32'b00001000011111011011111101010000;
		correct = 32'b01001001110011111011100010100101;
		#400 //1.2993701e-27 * 7.6359305e-34 = 1701652.6
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111110001000000001110100101;
		b = 32'b01000000001000110001011110101010;
		correct = 32'b10110111000110011101011010001010;
		#400 //-2.3366718e-05 * 2.5483193 = -9.169462e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001010001110010100110111101000;
		b = 32'b00010111011101111010010011010011;
		correct = 32'b00110010001111111000111010010110;
		#400 //8.9220785e-33 * 8.001804e-25 = 1.11500835e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100001111001010110101010000001;
		b = 32'b11101101111011110101101110011000;
		correct = 32'b10110011011101010101110111110100;
		#400 //5.2899735e+20 * -9.259706e+27 = -5.7128958e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111001111010001000111101011111;
		b = 32'b00101111110010001011000011101100;
		correct = 32'b11001001100101000101001101101101;
		#400 //-0.00044357308 * 3.65055e-10 = -1215085.6
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001111110111010011100000110101;
		b = 32'b01101010000000000111011011011001;
		correct = 32'b00100101010111000110101110001100;
		#400 //7422896600.0 * 3.8825937e+25 = 1.9118397e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011111100111101000111011001101;
		b = 32'b00110001110010011101111001011010;
		correct = 32'b11101101010010010001001101001101;
		#400 //-2.285059e+19 * 5.8751484e-09 = -3.8893638e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100000110101010001100101110101;
		b = 32'b01001111110011011110110110001010;
		correct = 32'b11010000100001000111010100101010;
		#400 //-1.2284346e+20 * 6909793300.0 = -17778168000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010110001010001111100110101000;
		b = 32'b11111101101011110011111110010110;
		correct = 32'b00010111111101101101011000010101;
		#400 //-46447555000000.0 * -2.9118132e+37 = 1.5951419e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100101111110100100000111011100;
		b = 32'b01000010011011111001101101101101;
		correct = 32'b01100011000001011011000001111011;
		#400 //1.4772581e+23 * 59.901783 = 2.4661337e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110000011001101111100010101;
		b = 32'b01000010101110011001011100010001;
		correct = 32'b00111010110000100101000011010110;
		#400 //0.13756974 * 92.79505 = 0.0014825116
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010001000010001100011011011101;
		b = 32'b01110111100000010111111101010101;
		correct = 32'b00011001000001110011000111111100;
		#400 //36715745000.0 * 5.253038e+33 = 6.989431e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000010100010100111001100110100;
		b = 32'b01010000101101111010000111101100;
		correct = 32'b10110001010000010000001011111000;
		#400 //-69.225006 * 24646738000.0 = -2.8086884e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011110001111101011010000001001;
		b = 32'b00001010001111011010011010100101;
		correct = 32'b01010011100000001011010111010001;
		#400 //1.0095747e-20 * 9.131361e-33 = 1105612400000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000100000110101000001011111110;
		b = 32'b10001011100011111101000000100000;
		correct = 32'b10111000000010011000010110110111;
		#400 //1.8162762e-36 * -5.539475e-32 = -3.2787877e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001110000100110001101111010001;
		b = 32'b11001101000011101101001011111000;
		correct = 32'b10000000100000111101011100000001;
		#400 //1.8132542e-30 * -149761920.0 = -1.2107579e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100111111011100100100001111011;
		b = 32'b01100011111111011010100110001000;
		correct = 32'b00000011011100000111101010101010;
		#400 //6.6136853e-15 * 9.3584845e+21 = 7.0670472e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111001001010101001100011001010;
		b = 32'b01011100010100100001101010011010;
		correct = 32'b00011100010011111101110011100001;
		#400 //0.00016269382 * 2.3655598e+17 = 6.8776034e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100001001101000101100011000011;
		b = 32'b00100101100001011111000110000111;
		correct = 32'b11111011001011000101100000011110;
		#400 //-2.0792562e+20 * 2.3235488e-16 = -8.948623e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011111110011110100011110110111;
		b = 32'b01011100011110101101110001010111;
		correct = 32'b11000010110100111000011011010000;
		#400 //-2.9872216e+19 * 2.8244404e+17 = -105.763306
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011011100001111110001001110000;
		b = 32'b01000110011111000110000100111000;
		correct = 32'b11010100100010011101010101101110;
		#400 //-7.6496185e+16 * 16152.305 = -4735930000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011100010000110101101001001000;
		b = 32'b10101111011001011100011001010010;
		correct = 32'b01101100010110011010011000110011;
		#400 //-2.1994754e+17 * -2.0897886e-10 = 1.052487e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000100011011111111001011110101;
		b = 32'b10000110011000110000100010001100;
		correct = 32'b01111101100001110100100000100010;
		#400 //-959.7962 * -4.2700234e-35 = 2.247754e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101001000011101010011111001000;
		b = 32'b00000010100111111001001001011111;
		correct = 32'b01100101111001001101110001110110;
		#400 //3.167586e-14 * 2.3446963e-37 = 1.3509579e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101010110001000001111110110011;
		b = 32'b10010001101010011100011011011110;
		correct = 32'b01011000100100111101110100100011;
		#400 //-3.483859e-13 * -2.678606e-28 = 1300623900000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101000000100010001011100110101;
		b = 32'b01100011000111111101011001111110;
		correct = 32'b10000100011010000110000101101011;
		#400 //-8.054149e-15 * 2.948488e+21 = -2.7316201e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101000111101111110101111000000;
		b = 32'b11001100100001000101001010111101;
		correct = 32'b11011011111011111101001000101010;
		#400 //9.366187e+24 * -69375464.0 = -1.35007195e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111100101110011000101001100001;
		b = 32'b11010111111111101010000110111010;
		correct = 32'b11100100001110101000100110011100;
		#400 //7.7070526e+36 * -559941130000000.0 = -1.3764041e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011100101100001110100111010011;
		b = 32'b10010011100100000100010110101110;
		correct = 32'b01001000100111001111010110101100;
		#400 //-1.1707145e-21 * -3.641942e-27 = 321453.38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101100101110000101001100110010;
		b = 32'b01001111011001010011101100111110;
		correct = 32'b10011100110011011101100101111111;
		#400 //-5.238831e-12 * 3845865000.0 = -1.3621983e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010110001001101111110010100010;
		b = 32'b00011010111011000001001111001100;
		correct = 32'b10111010101101010001010000110101;
		#400 //-1.348909e-25 * 9.7639296e-23 = -0.0013815226
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000001010111011010111111101000;
		b = 32'b10001010111011010000100111010000;
		correct = 32'b11110101111011110110101110111001;
		#400 //13.855446 * -2.2825961e-32 = -6.0700382e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001011001100010001011101110111;
		b = 32'b11011001011111010000111001000100;
		correct = 32'b10110001001100110010011011110000;
		#400 //11605879.0 * -4451803400000000.0 = -2.6070062e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101010110011001000010101000100;
		b = 32'b00110100010101010111110100000000;
		correct = 32'b10110101111101010011111100011110;
		#400 //-3.633015e-13 * 1.9882646e-07 = -1.8272292e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001010000111101011100010110101;
		b = 32'b10101111100111011101010100110000;
		correct = 32'b01011010000000001011100010000100;
		#400 //-2600493.2 * -2.8709612e-10 = 9057919000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100100101011111000011010110010;
		b = 32'b01000110011100111100111111111000;
		correct = 32'b00011101101110000100110011100001;
		#400 //7.6122335e-17 * 15603.992 = 4.8783885e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110010111101001000101110100100;
		b = 32'b11111111110000110001101111111001;
		correct = 32'b11111111110000110001101111111001;
		#400 //2.846884e-08 * nan = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011001100110111001011101110011;
		b = 32'b11011000010101011101000100111011;
		correct = 32'b11000000101110100100100110001101;
		#400 //5474392700000000.0 * -940378460000000.0 = -5.8214784
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100001011100011010101111101000;
		b = 32'b00000110111100011111010111001111;
		correct = 32'b11011001111111111011000111001111;
		#400 //-8.188149e-19 * 9.101531e-35 = -8996452700000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110110111110101100111110010;
		b = 32'b11001110010110001000101010001110;
		correct = 32'b00101000000001000000011010001010;
		#400 //-6.656389e-06 * -908239740.0 = 7.32889e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001110101011000010100101011101;
		b = 32'b11010001110101010101111001100000;
		correct = 32'b00111100010011101000111101001000;
		#400 //-1444196000.0 * -114551420000.0 = 0.012607403
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111000100000000001111110000010;
		b = 32'b11101100111100000000110110000101;
		correct = 32'b10001011000010001010001001110010;
		#400 //6.1093844e-05 * -2.3216483e+27 = -2.6314858e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000110100100110001101111101011;
		b = 32'b10011101011110011001111111101010;
		correct = 32'b10101000100101101101110110111110;
		#400 //5.5336276e-35 * -3.303755e-21 = -1.674951e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010010011101100111101101110001;
		b = 32'b00011110000000001011111101100110;
		correct = 32'b01110011111101010000110100000100;
		#400 //264658240000.0 * 6.815844e-21 = 3.8829856e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101100111000110110111110110111;
		b = 32'b01001110110111010101101011000011;
		correct = 32'b01011101100000111000010001010010;
		#400 //2.1996298e+27 * 1856856400.0 = 1.1845987e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011100101100100010100010001010;
		b = 32'b00000100111110101111101011101000;
		correct = 32'b01010111001101011011100011000011;
		#400 //1.1789531e-21 * 5.900514e-36 = 199805150000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010001011010011111010101001101;
		b = 32'b10011101110011110110110100101111;
		correct = 32'b10110011000100000101111101010010;
		#400 //1.8456048e-28 * -5.4905337e-21 = -3.3614306e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111011101001111101100111110100;
		b = 32'b10101111100111001100100101101100;
		correct = 32'b01001011100010010000100001110111;
		#400 //-0.0051224176 * -2.8519354e-10 = 17961198.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000110110100110111010001100;
		b = 32'b10111100110100000000101101101011;
		correct = 32'b00110011100001100110010000001001;
		#400 //-1.5893007e-09 * -0.02539607 = 6.2580575e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110110000101111111111101000101;
		b = 32'b11010011111101111111010010100111;
		correct = 32'b01100001100111001110110110100111;
		#400 //-7.707171e+32 * -2129923000000.0 = 3.618521e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100100011010010111100000010000;
		b = 32'b01100010100000010001001011101011;
		correct = 32'b11000001011001111000011011001010;
		#400 //-1.7226971e+22 * 1.1904966e+21 = -14.4704075
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101111100110111010010100111010;
		b = 32'b00000001001101111011011111100100;
		correct = 32'b11101101110110001110000111010101;
		#400 //-2.8311736e-10 * 3.3743727e-38 = -8.390222e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100100100010000100110111101010;
		b = 32'b10110010101111001100110000110001;
		correct = 32'b10110001001110001101001001100001;
		#400 //5.911259e-17 * -2.1978936e-08 = -2.689511e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110111000100010111100111101011;
		b = 32'b01110000100101000110101110011000;
		correct = 32'b11000101111110101110110000001001;
		#400 //-2.9506087e+33 * 3.6747083e+29 = -8029.5044
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100001111000000011010101010110;
		b = 32'b01001011011001111100010101111110;
		correct = 32'b10010101111101111010010101110010;
		#400 //-1.5192948e-18 * 15189374.0 = -1.0002353e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000100011010001111000001001101;
		b = 32'b00000001100000111010011111001111;
		correct = 32'b01000010011000100111100010010010;
		#400 //2.738181e-36 * 4.8362594e-38 = 56.617744
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100101111011110000111110011011;
		b = 32'b00100010011010110000011101010011;
		correct = 32'b11000011000000100011001000110010;
		#400 //-4.1470466e-16 * 3.1852316e-18 = -130.19608
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001111001101100100001010000010;
		b = 32'b10011100001010100101001101011111;
		correct = 32'b11110010100010001111011111110001;
		#400 //3057812000.0 * -5.6356036e-22 = -5.425882e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001010011000011101011110110111;
		b = 32'b01011000110001011100111101000101;
		correct = 32'b00110001000100100010001111001000;
		#400 //3700205.8 * 1739952000000000.0 = 2.1266136e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001010100110010010011000011100;
		b = 32'b01100101111010010000011101011000;
		correct = 32'b00100100001010000011111011110000;
		#400 //5018382.0 * 1.3755586e+23 = 3.6482503e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010001010111101011101101001;
		b = 32'b10011111001111001101111111100001;
		correct = 32'b01011010011010001110100111010101;
		#400 //-0.0006555231 * -3.9995737e-20 = 1.6389824e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011111000001100111100101110;
		b = 32'b10110011011110001101001000011011;
		correct = 32'b01010111111001110100101110110111;
		#400 //-29466204.0 * -5.793309e-08 = 508624760000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010001101101110011110001111101;
		b = 32'b10010010011011001100010101101001;
		correct = 32'b00111110110001100001111000010000;
		#400 //-2.8909588e-28 * -7.4711796e-28 = 0.3869481
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011101111000110010010111101000;
		b = 32'b01010100100011100000001100101111;
		correct = 32'b00001000110011001011110000111010;
		#400 //6.0125594e-21 * 4879510000000.0 = 1.2322055e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110010000100010000000101101001;
		b = 32'b01001100111011000000101110010010;
		correct = 32'b01100100100111010100001110010101;
		#400 //2.87213e+30 * 123755660.0 = 2.320807e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110000000111100011010111101000;
		b = 32'b01111110111011000110010101101101;
		correct = 32'b00110000101010110101010010100011;
		#400 //1.958552e+29 * 1.5711222e+38 = 1.2465943e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000000100010001111001100011010;
		b = 32'b11100011011111111101000110111011;
		correct = 32'b00011100100010010000101111011111;
		#400 //-4.2796755 * -4.7190324e+21 = 9.068968e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100110110111011110110001111111;
		b = 32'b01101000001011000101011111100001;
		correct = 32'b00111110001001001101001011011011;
		#400 //5.240028e+23 * 3.2554725e+24 = 0.1609606
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101111111000001010001101001011;
		b = 32'b10111001011100001100010001011101;
		correct = 32'b11110101111011101101100110110001;
		#400 //1.390441e+29 * -0.00022961335 = -6.055576e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010111111100111110111111011100;
		b = 32'b01000001010010100000110011110010;
		correct = 32'b10010110000110101000100100000100;
		#400 //-1.5764056e-24 * 12.62816 = -1.2483255e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111100111101001001000101101000;
		b = 32'b00101001001010101110110000011000;
		correct = 32'b11010011001101110010011011010111;
		#400 //-0.029854491 * 3.795236e-14 = -786630640000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000110101110101000011101101010;
		b = 32'b00111011100001110100101111001101;
		correct = 32'b11001010101100000111100001010100;
		#400 //-23875.707 * 0.004128909 = -5782570.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001000111011111000010100110000;
		b = 32'b00110110111110011110000000000100;
		correct = 32'b10010001011101010110010000110010;
		#400 //-1.44156015e-33 * 7.446857e-06 = -1.9357967e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100001011010110001011010111000;
		b = 32'b01001100011101110101110110101010;
		correct = 32'b11010100011100110100101101011010;
		#400 //-2.7103887e+20 * 64845480.0 = -4179765000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001001110110010101000011011001;
		b = 32'b11111111000101101011100001100001;
		correct = 32'b00001010001110001000111010000010;
		#400 //-1780251.1 * -2.0034155e+38 = 8.8860805e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110010001000000011011111010110;
		b = 32'b10101001010101101011010011101110;
		correct = 32'b11001000001111110000100000101001;
		#400 //9.325921e-09 * -4.7674477e-14 = -195616.64
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010101100000110110101011001001;
		b = 32'b01000110111010000011011000110101;
		correct = 32'b01001110000100001110000100111001;
		#400 //18061833000000.0 * 29723.104 = 607669800.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111110100001110001000101010100;
		b = 32'b11100100101101101100011010101100;
		correct = 32'b00011001001111010010110110111100;
		#400 //-0.26380408 * -2.6972986e+22 = 9.780307e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110010011010011001011100110011;
		b = 32'b10000000010110000110000111101111;
		correct = 32'b01110001101010010010011000010110;
		#400 //-1.3596764e-08 * -8.116656e-39 = 1.6751683e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110011100000110000101111000111;
		b = 32'b10100011010101011110110101010110;
		correct = 32'b11001111100111001101000110011001;
		#400 //6.102305e-08 * -1.1597011e-17 = -5261964000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110011100100010000000100000010;
		b = 32'b01011101000110110001000010110111;
		correct = 32'b10010101111011110110001110111000;
		#400 //-6.752272e-08 * 6.98352e+17 = -9.668866e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011110000111001010001101100100;
		b = 32'b10001100110100001011101010100101;
		correct = 32'b11010000110000000001110010110101;
		#400 //8.29236e-21 * -3.2159807e-31 = -25784855000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010000111011000101110011101101;
		b = 32'b00101010101011011111110110111101;
		correct = 32'b01100101101011011110001010010011;
		#400 //31724104000.0 * 3.090704e-13 = 1.0264362e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111111101010001111111001101001;
		b = 32'b11110001101000111000100010011100;
		correct = 32'b10001101100001000100011000010100;
		#400 //1.320264 * -1.6195586e+30 = -8.151999e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001100000100000110001011101110;
		b = 32'b10011001011111001110101110010101;
		correct = 32'b01110010000100100010010100000101;
		#400 //-37850040.0 * -1.307567e-23 = 2.8946922e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101100100010100110101010111011;
		b = 32'b00000111100011010001010011111011;
		correct = 32'b11100100011110110010101000000110;
		#400 //-3.9340454e-12 * 2.1227653e-34 = -1.8532643e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100110111111010110001001100100;
		b = 32'b10111011111101001001000010101011;
		correct = 32'b00101010100001001001110110100100;
		#400 //-1.758207e-15 * -0.007463535 = 2.3557295e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100011111000000011001001011110;
		b = 32'b10110000001111101000001101001111;
		correct = 32'b10110011000101101010000110010100;
		#400 //2.430746e-17 * -6.93082e-10 = -3.507155e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101000011100011011100010000011;
		b = 32'b00101101010100101101110100011001;
		correct = 32'b00111010100100101011101100101001;
		#400 //1.3418197e-14 * 1.19862115e-11 = 0.0011194694
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010100001000110110001010011111;
		b = 32'b10111001100000100111100100011111;
		correct = 32'b01011010001000000100100111001011;
		#400 //-2806937000000.0 * -0.00024885774 = 1.1279283e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011101001010011110110110010000;
		b = 32'b10101010111000111001100101011110;
		correct = 32'b00110001101111110010000111100110;
		#400 //-2.248978e-21 * -4.042972e-13 = 5.5626854e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101110111010100100101000011100;
		b = 32'b10000101000010001101110000100111;
		correct = 32'b11101001010110110001111101000111;
		#400 //1.06542525e-10 * -6.435125e-36 = -1.6556404e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100001110111011011110111010000;
		b = 32'b00101010110101101100101011000000;
		correct = 32'b10110110100001000010010000110000;
		#400 //-1.5025785e-18 * 3.8154722e-13 = -3.9381193e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101001011011110000001101110111;
		b = 32'b10101011100000000011000110101001;
		correct = 32'b00111101011011101010011011100000;
		#400 //-5.3071666e-14 * -9.10873e-13 = 0.058264613
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010101010001101111000111110011;
		b = 32'b10011001101010110010010101100101;
		correct = 32'b01111011000101001100101001110111;
		#400 //-13671404000000.0 * -1.7696089e-23 = 7.725664e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100110011001100101001111011001;
		b = 32'b01001110100101001000000101000110;
		correct = 32'b11010111010001101000011001011011;
		#400 //-2.7192275e+23 * 1245750000.0 = -218280350000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000100111001010111011110000001;
		b = 32'b00011000101111100001001011010001;
		correct = 32'b10101011100110101000011101000100;
		#400 //-5.394739e-36 * 4.913285e-24 = -1.0979902e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111110000111010101001100010;
		b = 32'b10100001011000000000001100010011;
		correct = 32'b11100101110111111001101100010101;
		#400 //100180.766 * -7.589822e-19 = -1.3199356e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001111001100111110110001101101;
		b = 32'b10000011100111000111010001011011;
		correct = 32'b11001011000100110011001101100001;
		#400 //8.870915e-30 * -9.19557e-37 = -9646945.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011101110101011000010001010001;
		b = 32'b01001000110011011010001100011111;
		correct = 32'b10010100100001001110011110011101;
		#400 //-5.6517443e-21 * 421144.97 = -1.3419949e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011111111111010111100111010000;
		b = 32'b00001011110100100000110101000110;
		correct = 32'b01010011100110100111011000011111;
		#400 //1.0735119e-19 * 8.090903e-32 = 1326813400000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001100011001000000001111101010;
		b = 32'b11101011011000001001110000100000;
		correct = 32'b10100000100000011111000011010000;
		#400 //59772840.0 * -2.7153666e+26 = -2.2012806e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100101101000100010010101110110;
		b = 32'b10001011001010000100110111110110;
		correct = 32'b11011001111101101010001000010000;
		#400 //2.8127905e-16 * -3.2414274e-32 = -8677629000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000111011111011110010010010010;
		b = 32'b00010011110001111010101000110101;
		correct = 32'b11110011001000101100001110100000;
		#400 //-64996.57 * 5.04025e-27 = -1.2895505e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000100011111001111010000100011;
		b = 32'b11000010111111010001000011101100;
		correct = 32'b00000000111111111110001011100010;
		#400 //-2.973456e-36 * -126.53305 = 2.3499442e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110010101001111001010010110010;
		b = 32'b01110111011011111001001010000111;
		correct = 32'b10111010101100110001001001101100;
		#400 //-6.638561e+30 * 4.859105e+33 = -0.0013662106
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101110011000000000100000000000;
		b = 32'b11001001100100101010000010110011;
		correct = 32'b10100100010000111001000111110010;
		#400 //5.093881e-11 * -1201174.4 = -4.2407505e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101110100100001000000111011110;
		b = 32'b01000001000110001011110101001101;
		correct = 32'b00101100111100100011001111010010;
		#400 //6.571431e-11 * 9.546216 = 6.883807e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001110101011000001010110001001;
		b = 32'b00001000011001111110011001111110;
		correct = 32'b11000101101111011111011110101111;
		#400 //-4.242201e-30 * 6.9784976e-34 = -6078.9604
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001110111100011010110001100011;
		b = 32'b10111010100111001010100100011010;
		correct = 32'b11010011110001010111010111000011;
		#400 //2027303300.0 * -0.0011952252 = -1696168500000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110101101110110001000000101100;
		b = 32'b10011100111100101001100110101111;
		correct = 32'b11011000010001010110010100110100;
		#400 //1.3937292e-06 * -1.6053943e-21 = -868153800000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010010111101101110001011110000;
		b = 32'b11100000101000001101000110000001;
		correct = 32'b10110001110001001000000100001100;
		#400 //530184670000.0 * -9.270548e+19 = -5.7190217e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111000011001011100010011011100;
		b = 32'b11011100001100101000000001101101;
		correct = 32'b10011011101001001100001101000101;
		#400 //5.4781194e-05 * -2.00975e+17 = -2.7257714e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110111001110000011101010001011;
		b = 32'b10011111101111011111001101110110;
		correct = 32'b11010110111110000100100110110101;
		#400 //1.0980885e-05 * -8.0447386e-20 = -136497730000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101111101001101111100101011001;
		b = 32'b11111101110100110100010101101010;
		correct = 32'b00110001010010100101001100011000;
		#400 //-1.0335191e+29 * -3.510344e+37 = 2.9442102e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001011100010001111110101110000;
		b = 32'b00000010000010010000000111110100;
		correct = 32'b01001000111111111111011110010000;
		#400 //5.2766625e-32 * 1.0065731e-37 = 524220.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101000111110010010011011010100;
		b = 32'b01100100111100100001100100110110;
		correct = 32'b10000011100000111011101010100110;
		#400 //-2.7661392e-14 * 3.572743e+22 = -7.74234e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101001000101011011111111000101;
		b = 32'b10000111001000010110001101101010;
		correct = 32'b11100001011011011000100110010101;
		#400 //3.325098e-14 * -1.2141509e-34 = -2.7386201e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101100001010110000011001111000;
		b = 32'b00111111101010000111100011011110;
		correct = 32'b11101100000000011111000010010110;
		#400 //-8.2702745e+26 * 1.3161886 = -6.2835026e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100001101100110101101001100100;
		b = 32'b11111111110100101000100100011111;
		correct = 32'b11111111110100101000100100011111;
		#400 //-4.1356007e+20 * nan = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110100101110011011110000011;
		b = 32'b00011111001100001111011000011111;
		correct = 32'b11010110110110101100000110111110;
		#400 //-4.506613e-06 * 3.7473036e-20 = -120262826000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001000110001001111000011101111;
		b = 32'b10111101100111110000110110110010;
		correct = 32'b11001010100111100111110110010001;
		#400 //403335.47 * -0.07766284 = -5193416.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001100111011110110001101110010;
		b = 32'b00110101001110000001000011000100;
		correct = 32'b11010111001001100111100011001011;
		#400 //-125508500.0 * 6.856974e-07 = -183037730000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100000101011110010101001010000;
		b = 32'b01011011111101100100111011001001;
		correct = 32'b01000100001101100000111011011101;
		#400 //1.0097591e+20 * 1.3865894e+17 = 728.23224
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010111010001111000000110100;
		b = 32'b00111000101001011110010011011100;
		correct = 32'b11000001101100111011101011011000;
		#400 //-0.0017771781 * 7.9104415e-05 = -22.466232
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101010110101111001111001101111;
		b = 32'b10110110001011110100011101000101;
		correct = 32'b10110100000111010111010110010110;
		#400 //3.8301607e-13 * -2.6118516e-06 = -1.4664542e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111001110110001101100001110101;
		b = 32'b11110111000101000000010001101011;
		correct = 32'b00000010001110111000010100101101;
		#400 //-0.00041360004 * -3.0021466e+33 = 1.377681e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110011001001110010011000011111;
		b = 32'b01010110000100011011100100010111;
		correct = 32'b01011100100100101101000111101111;
		#400 //1.3242901e+31 * 40056035000000.0 = 3.3060937e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110001010010100110111100100000;
		b = 32'b11100110100101000110100000101100;
		correct = 32'b01001010001011101001100100011011;
		#400 //-1.002405e+30 * -3.5041594e+23 = 2860614.8
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111111011101110011111010001001;
		b = 32'b11111001000100001111111000011000;
		correct = 32'b01000101110110100100010010101011;
		#400 //-3.2864402e+38 * -4.7052774e+34 = 6984.5835
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001101011111010000011001010111;
		b = 32'b01000011011100101001010001010111;
		correct = 32'b10001001100001011000001011111000;
		#400 //-7.7969275e-31 * 242.57945 = -3.2141748e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101111000001111011100010010000;
		b = 32'b01101110011011010101111010111100;
		correct = 32'b11000000000100100101111101111100;
		#400 //-4.20036e+28 * 1.8365619e+28 = -2.287078
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111110001011100111001000111110;
		b = 32'b00101001110010101100011100100001;
		correct = 32'b11010011110111000011101101111011;
		#400 //-0.17035767 * 9.0051454e-14 = -1891781400000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101100110011000100011001000001;
		b = 32'b11111000101001110001111101101101;
		correct = 32'b10110011100111000111010001100010;
		#400 //1.975621e+27 * -2.7117218e+34 = -7.285486e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110100111010011100111110111111;
		b = 32'b00010100101011111000000010110101;
		correct = 32'b11011111101010101000011011001001;
		#400 //-4.3550787e-07 * 1.772125e-26 = -2.457546e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110101010100101101101011001;
		b = 32'b00110111001100011111100000110000;
		correct = 32'b10111110111101010000110010110010;
		#400 //-5.077029e-06 * 1.0607808e-05 = -0.47861248
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011001011001110010110101100000;
		b = 32'b11111010001001000011011110011001;
		correct = 32'b00011110101101000011000101000001;
		#400 //-4066913000000000.0 * -2.1316608e+35 = 1.9078612e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100010001110100110110111000010;
		b = 32'b01011110010111011101011010000101;
		correct = 32'b10000011010101110010001101001110;
		#400 //-2.5265806e-18 * 3.9962775e+18 = -6.322335e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010101011110011010110100111000;
		b = 32'b10110111011101110000010000100000;
		correct = 32'b01011101100000010110000011101111;
		#400 //-17157648000000.0 * -1.4723308e-05 = 1.1653393e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110101001001000101011101101110;
		b = 32'b10110011111001000010100000000000;
		correct = 32'b01000000101110000110010110111111;
		#400 //-6.122199e-07 * -1.0624353e-07 = 5.76242
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101110011100101000110111101100;
		b = 32'b01010100001111010010100111011010;
		correct = 32'b00011001101001000010000010101111;
		#400 //5.515048e-11 * 3249804000000.0 = 1.6970403e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101101000100110010101001000100;
		b = 32'b01100010111011000001110010101101;
		correct = 32'b10001001100111111000111110011101;
		#400 //-8.365367e-12 * 2.177749e+21 = -3.841291e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011110010000101001001101001110;
		b = 32'b10010000111100000001011111010011;
		correct = 32'b11001100110011110111011101110111;
		#400 //1.0300736e-20 * -9.4700016e-29 = -108772280.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000101110001000100000011001000;
		b = 32'b10111010110011010101010011100000;
		correct = 32'b01001010011101001010111001100111;
		#400 //-6280.0977 * -0.0015665554 = 4008857.8
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110101000010000000101100000101;
		b = 32'b01110011001110001101101010101111;
		correct = 32'b01000001001111000110011100010001;
		#400 //1.7245505e+32 * 1.4645661e+31 = 11.775163
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000000011011111001110100000110;
		b = 32'b10100001010010100010100011010111;
		correct = 32'b10011110100011010101011011001000;
		#400 //1.025007e-38 * -6.8494313e-19 = -1.4964848e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011000101101101000101000000001;
		b = 32'b10011111110011011001110111110111;
		correct = 32'b10111000011000110100010001100101;
		#400 //4.7185246e-24 * -8.708221e-20 = -5.4184715e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010111101110110101111101000111;
		b = 32'b00011011011000001100110100111001;
		correct = 32'b11111011110101010110000001000010;
		#400 //-412035770000000.0 * 1.8595157e-22 = -2.2158231e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001010101110111010000110000101;
		b = 32'b01000000111010101101001001101110;
		correct = 32'b01001001010011001000110110001011;
		#400 //6148290.5 * 7.338187 = 837848.7
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000111000111010011000001000111;
		b = 32'b01000000111000011001001110011110;
		correct = 32'b10000101101100100110001101110101;
		#400 //-1.1825555e-34 * 7.0492697 = -1.6775574e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100010001101110011000000000111;
		b = 32'b10001100100000111101010101111111;
		correct = 32'b11010101001100011101110000110101;
		#400 //2.482655e-18 * -2.031224e-31 = -12222459000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101001011011010010100000100011;
		b = 32'b10110110111100000101011101010100;
		correct = 32'b10110001111111001001101110110010;
		#400 //5.2659384e-14 * -7.1627237e-06 = -7.351866e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011010101011000110111011011000;
		b = 32'b10110001100010001110010001000000;
		correct = 32'b00101000101000010011101110011011;
		#400 //-7.131661e-23 * -3.98407e-09 = 1.790044e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000011000001111011000001100100;
		b = 32'b11110010100100110001101001000010;
		correct = 32'b00001111111011000010001100100000;
		#400 //-135.68903 * -5.827333e+30 = 2.3284926e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101010110011101111011100111010;
		b = 32'b11011010011100100110000010011111;
		correct = 32'b01001111110110101001100100011000;
		#400 //-1.2510311e+26 * -1.7055795e+16 = 7334932500.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010001010111101011010010111010;
		b = 32'b01010100110001110111101111011111;
		correct = 32'b10111100000011101110011010001101;
		#400 //-59782177000.0 * 6854213600000.0 = -0.00872196
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000101010101011111010110001111;
		b = 32'b00000100100001011011010000101001;
		correct = 32'b01000000010011001101010011110001;
		#400 //1.0060314e-35 * 3.14336e-36 = 3.200497
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101001010111011110001110101111;
		b = 32'b01101000110010011001000110100111;
		correct = 32'b01000000000011001110011101100011;
		#400 //1.6765488e+25 * 7.61506e+24 = 2.2016227
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100101101001000101111001011111;
		b = 32'b01000100100011001010000100100001;
		correct = 32'b10100000100101011001101101111000;
		#400 //-2.8513413e-16 * 1125.0353 = -2.5344462e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001111110111010001001011111000;
		b = 32'b00010000100000000011001000110110;
		correct = 32'b01111110110111001011110001100001;
		#400 //7418016000.0 * 5.056446e-29 = 1.4670414e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110011111111011110111000110011;
		b = 32'b11001111010110101100011101011010;
		correct = 32'b10100100000101001001000011101100;
		#400 //1.1824559e-07 * -3670497800.0 = -3.2215138e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001110010101101110100011101110;
		b = 32'b11000101010000000000000010111101;
		correct = 32'b00001000100011110100010101100111;
		#400 //-2.6489688e-30 * -3072.0461 = 8.622816e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110001110110010010010001010110;
		b = 32'b00110110010111101101010011101110;
		correct = 32'b11111010111110010111011010011000;
		#400 //-2.1504696e+30 * 3.320452e-06 = -6.4764364e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111001101010010111111011011101;
		b = 32'b01010100010100000000111101110101;
		correct = 32'b00100100110100001000110010100100;
		#400 //0.00032328712 * 3574450000000.0 = 9.0443875e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101101111111000010100101010001;
		b = 32'b10010011011110010001100110111011;
		correct = 32'b11011010000000011001001010100101;
		#400 //2.8667431e-11 * -3.1440905e-27 = -9117877000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100100111111100011111110110000;
		b = 32'b11011100110110010111001111110101;
		correct = 32'b01000111100101011010100011000100;
		#400 //-3.7520497e+22 * -4.8966053e+17 = 76625.53
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010000111100000101001011010100;
		b = 32'b01110101100010000011110110101111;
		correct = 32'b00011010111000011100100101101110;
		#400 //32255680000.0 * 3.4541185e+32 = 9.3383246e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101101001111011001011101111010;
		b = 32'b11100111010011010010100000110010;
		correct = 32'b00000101011011001001001111000101;
		#400 //-1.0777041e-11 * -9.688266e+23 = 1.1123808e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111011101001001000011010000001;
		b = 32'b11100101111000001011001111110100;
		correct = 32'b00010101001110110111000011011010;
		#400 //-0.005020917 * -1.32641205e+23 = 3.7853373e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001001101110100000000001111100;
		b = 32'b11011001100001111001000011111100;
		correct = 32'b10101111101011111001111011011111;
		#400 //1523727.5 * -4769817000000000.0 = -3.19452e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001101001101011001011001000110;
		b = 32'b10111011101000010010010111000011;
		correct = 32'b11010001000100000011110000110100;
		#400 //190407780.0 * -0.0049178316 = -38717833000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111100000010111011010011000000;
		b = 32'b01010101001100000000001101001111;
		correct = 32'b11100110010010110011000110100010;
		#400 //-2.9015812e+36 * 12095516000000.0 = -2.3988899e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111001101001010010000001001101;
		b = 32'b01111111011010100100000111000100;
		correct = 32'b00111001101101000111001111100111;
		#400 //1.0717301e+35 * 3.1138083e+38 = 0.0003441863
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000010100110101110000000001101;
		b = 32'b01011010100101001100000101001000;
		correct = 32'b10100111100001010100010000101011;
		#400 //-77.4376 * 2.0935406e+16 = -3.6988823e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011100001111111001001100101;
		b = 32'b11011010000111000100000001111101;
		correct = 32'b00110000110111101011101110001100;
		#400 //-17818826.0 * -1.099525e+16 = 1.620593e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001110001010111111100011001011;
		b = 32'b10100010001110101100100011101100;
		correct = 32'b01101011011010111011001010101000;
		#400 //-721302200.0 * -2.5314068e-18 = 2.8494125e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010111010111000110111101100000;
		b = 32'b10110101111110111000101010001111;
		correct = 32'b01100000111000000101011110101010;
		#400 //-242370910000000.0 * -1.8741283e-06 = 1.2932461e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010100101001100011000101110000;
		b = 32'b10101110100001100110000111111101;
		correct = 32'b01100101100111100100110010101001;
		#400 //-5710352000000.0 * -6.111021e-11 = 9.34435e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101100110011101000110011001001;
		b = 32'b11011110110111111100111111001000;
		correct = 32'b01001101011011000100000101111000;
		#400 //-1.9976285e+27 * -8.0636643e+18 = 247732100.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001100011100000000101100011100;
		b = 32'b00101010101110010010001111110100;
		correct = 32'b00100001001001011111010101000110;
		#400 //1.849227e-31 * 3.288755e-13 = 5.622879e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000011001001101010001101000010;
		b = 32'b10001101011110110010111001101110;
		correct = 32'b01110101001010011101010110100001;
		#400 //-166.63773 * -7.7401234e-31 = 2.152908e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100011011101101110110110001110;
		b = 32'b01011101001100100101100001111000;
		correct = 32'b00000101101100010011100011011011;
		#400 //1.3385991e-17 * 8.031971e+17 = 1.6665885e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011101101010010001101111011000;
		b = 32'b01110001010111111110011110011110;
		correct = 32'b10101011110000010101100101110000;
		#400 //-1.5231963e+18 * 1.10872264e+30 = -1.3738299e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010011111011110001110101101010;
		b = 32'b11110110000100001000101011111010;
		correct = 32'b10011101010100111011111110010000;
		#400 //2053981300000.0 * -7.3291946e+32 = -2.8024653e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101000110100001011001010001110;
		b = 32'b10110110011110010101000100010001;
		correct = 32'b01110001110101100100101010111101;
		#400 //-7.884368e+24 * -3.7151078e-06 = 2.1222446e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011011010001010111010111111111;
		b = 32'b01000110110011000000000011000110;
		correct = 32'b00010011111101111100101001011010;
		#400 //1.6333585e-22 * 26112.387 = 6.25511e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001011110111101110101000010000;
		b = 32'b10110110110111010001011011101101;
		correct = 32'b11010100100000010000111001110011;
		#400 //29217824.0 * -6.588982e-06 = -4434345600000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111100001010110010000010100011;
		b = 32'b01101110100101110001010001000110;
		correct = 32'b11001101000100001111110001010101;
		#400 //-3.554179e+36 * 2.3378373e+28 = -152028500.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100111110010011111110011100000;
		b = 32'b11001011001011110111111000110010;
		correct = 32'b10011100000100110101001100011100;
		#400 //5.6062875e-15 * -11501106.0 = -4.8745636e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011111011010000000011011101001;
		b = 32'b10111001001011110001010011110000;
		correct = 32'b11100101101010011010000111000100;
		#400 //1.6719307e+19 * -0.000166971 = -1.00133e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101000011101011001110100100100;
		b = 32'b11011111110010111000101000100010;
		correct = 32'b00001000000110100111010110010001;
		#400 //-1.36343065e-14 * -2.9333145e+19 = 4.648089e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001110001001001011001100011111;
		b = 32'b10110001011111101001100010110010;
		correct = 32'b00011100001001011001101110001111;
		#400 //-2.0300804e-30 * -3.7048662e-09 = 5.4794975e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110100110011110010101011001010;
		b = 32'b11101001110011000110011011111111;
		correct = 32'b00001010100000011011101100111011;
		#400 //-3.8587888e-07 * -3.0888407e+25 = 1.2492676e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001010111110011100001010111110;
		b = 32'b11000010001101100111111110011010;
		correct = 32'b11001000001011110010110100010111;
		#400 //8184159.0 * -45.62461 = -179380.36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010111010001101111111000001111;
		b = 32'b01001111100101111000011111100001;
		correct = 32'b10000111001010000001011101101010;
		#400 //-6.4297918e-25 * 5084529000.0 = -1.2645796e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000001010011110000111010011101;
		b = 32'b01111100110011000110110100001111;
		correct = 32'b10000100000000011010010110111110;
		#400 //-12.941068 * 8.491524e+36 = -1.5239982e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010011101100001100010100010100;
		b = 32'b10011010011101001001001001111100;
		correct = 32'b10111000101110010000011110001111;
		#400 //4.462298e-27 * -5.0576347e-23 = -8.822895e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110011101000011010011000111010;
		b = 32'b11100111100111111000111001101010;
		correct = 32'b00001011100000011010110111011000;
		#400 //-7.527383e-08 * -1.5069667e+24 = 4.9950564e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100100100100000001101001100001;
		b = 32'b01011110110011101000010110000110;
		correct = 32'b00000101001100101010000010010011;
		#400 //6.249473e-17 * 7.440724e+18 = 8.3990126e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000110111111111000100111011111;
		b = 32'b10010101111110111110010110100010;
		correct = 32'b00110000100000011101100110110110;
		#400 //-9.612292e-35 * -1.0174039e-25 = 9.447862e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111001100001101111101010011110;
		b = 32'b11010111100000011100101001001011;
		correct = 32'b01100001100001010001111000000001;
		#400 //-8.760636e+34 * -285411700000000.0 = 3.0694737e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010011100110111111000000001000;
		b = 32'b01000100101110111011110000010111;
		correct = 32'b10001110010101001010010000000001;
		#400 //-3.936419e-27 * 1501.8778 = -2.6209982e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001000110111000000010000101110;
		b = 32'b00000100011010111000100011110110;
		correct = 32'b01000011111011110010001000001001;
		#400 //1.3241751e-33 * 2.7687007e-36 = 478.2659
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011001011011111011111110011101;
		b = 32'b01011110111111000101111001010101;
		correct = 32'b00111001111100110011001011001011;
		#400 //4217700000000000.0 * 9.092533e+18 = 0.00046386415
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001001001010011110100000011110;
		b = 32'b10101101101110101011110010011100;
		correct = 32'b01011010111010001110110101101110;
		#400 //-695937.9 * -2.1229511e-11 = 3.2781626e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110010000001101110110010011011;
		b = 32'b10010101001110110011000100011011;
		correct = 32'b11011100001110001000010100010101;
		#400 //7.853624e-09 * -3.7803087e-26 = -2.0775088e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111101001111010001111000100;
		b = 32'b00101001100111101101010100111111;
		correct = 32'b11001101100001110001100011011110;
		#400 //-1.998421e-05 * 7.053602e-14 = -283319230.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100001111010110101001000010111;
		b = 32'b11101010101000110110001000100001;
		correct = 32'b10110110101110000101101110101111;
		#400 //5.426125e+20 * -9.8759155e+25 = -5.4943007e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011101100011001111111100001011;
		b = 32'b11001110000011110101101110000010;
		correct = 32'b01001110111110111100100010010100;
		#400 //-1.2699814e+18 * -601284740.0 = 2112113200.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000100110001110011010000010110;
		b = 32'b10111011011100111110001110000010;
		correct = 32'b01001000110100010001100010000010;
		#400 //-1593.6277 * -0.0037214463 = 428228.06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001100000000010101000011100010;
		b = 32'b11000000011011000000010010100110;
		correct = 32'b11001011000011000100001110011110;
		#400 //33899400.0 * -3.6877837 = -9192350.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110010101110100111100010101011;
		b = 32'b10110111001000011011010111110101;
		correct = 32'b00111011000100111001100101010010;
		#400 //-2.1708123e-08 * -9.638713e-06 = 0.0022521806
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111100101010001001001010111111;
		b = 32'b11111111111010111000111001100011;
		correct = 32'b11111111111010111000111001100011;
		#400 //-7.002258e+36 * nan = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101001010110101111010110101011;
		b = 32'b10110101001010111110000101111111;
		correct = 32'b10110011101000110000111101000111;
		#400 //4.8618807e-14 * -6.4030604e-07 = -7.593058e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111010101100000111001010100000;
		b = 32'b11111011000100101000111010000111;
		correct = 32'b10111111000110100001101100110100;
		#400 //4.5808456e+35 * -7.609661e+35 = -0.6019776
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010100100101000111011011111010;
		b = 32'b00111111101101001011010100011001;
		correct = 32'b00010100010100100101001011000011;
		#400 //1.4991109e-26 * 1.4117767 = 1.06186124e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110001110111100111010101101001;
		b = 32'b01010111111111011110001110101111;
		correct = 32'b11011001011000000100111011010110;
		#400 //-2.2031236e+30 * 558308670000000.0 = -3946067200000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000101110100010000101001001111;
		b = 32'b00101001001111111101011101110110;
		correct = 32'b01011100000010110111100110101000;
		#400 //6689.2886 * 4.2597402e-14 = 1.5703514e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001010101100111111011101011010;
		b = 32'b10111101100000111011100111000111;
		correct = 32'b00001100101011101110000001001000;
		#400 //-1.7330116e-32 * -0.064319186 = 2.694393e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011101010110010000001010101000;
		b = 32'b01101000110100000001010111001010;
		correct = 32'b00110100000001010111110101111111;
		#400 //9.7732785e+17 * 7.8612333e+24 = 1.2432245e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010100001100110010011000011101;
		b = 32'b11101001111010010001011101110011;
		correct = 32'b00101001110001001100000101111001;
		#400 //-3077754300000.0 * -3.5223806e+25 = 8.737711e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110000111101010111000010110001;
		b = 32'b00101011010010001111110001011001;
		correct = 32'b01000101000111000100111110110011;
		#400 //1.7858125e-09 * 7.1404476e-13 = 2500.9812
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100010001010100110011001000001;
		b = 32'b01010111110110001101001011011001;
		correct = 32'b00001001110010010011000000001111;
		#400 //2.3093429e-18 * 476800200000000.0 = 4.8434184e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100101000010110100110100010010;
		b = 32'b01001100100001101011110101111010;
		correct = 32'b10011000000001000101010100110000;
		#400 //-1.208244e-16 * 70642640.0 = -1.7103609e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101001111011101010010100110101;
		b = 32'b11111110000101010101011010011110;
		correct = 32'b00101011010011001000101111011001;
		#400 //-3.6063064e+25 * -4.962618e+37 = 7.2669437e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110011110001101001011100110100;
		b = 32'b01100100010000110110011101010100;
		correct = 32'b10001111000000100001011001110001;
		#400 //-9.247597e-08 * 1.4418243e+22 = -6.413817e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000111000111110001100101100101;
		b = 32'b10100100000110010101010100010100;
		correct = 32'b00100010100001001101000001101001;
		#400 //-1.1969293e-34 * -3.324865e-17 = 3.5999335e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111110011011010100000010111011;
		b = 32'b11011100000011100110110111110100;
		correct = 32'b11100001110101010011011110000001;
		#400 //7.8840784e+37 * -1.6036137e+17 = -4.916445e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001010111101101011001101101110;
		b = 32'b01100011111010011101100111110110;
		correct = 32'b00100110100001110000100010000011;
		#400 //8083895.0 * 8.627594e+21 = 9.369814e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011000100000110010101010111;
		b = 32'b10110010100101100111000010011000;
		correct = 32'b01010111111101011011011100010011;
		#400 //-9463127.0 * -1.75135e-08 = 540333300000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000011110100001011000010001000;
		b = 32'b01000101101110111110001110000100;
		correct = 32'b10111101100011100010101110110001;
		#400 //-417.37915 * 6012.4395 = -0.06941927
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000010010101000001010110111011;
		b = 32'b00101101101011111010101001001100;
		correct = 32'b00010100000110101000100110011010;
		#400 //1.5581536e-37 * 1.9970824e-11 = 7.80215e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100100010100011111001010100100;
		b = 32'b01111010011010001010001110100000;
		correct = 32'b10101001011001110000011110110010;
		#400 //-1.5491414e+22 * 3.019829e+35 = -5.129898e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001000001011110100101110000001;
		b = 32'b00100100000101110111011110111000;
		correct = 32'b11100011100101000010001010110111;
		#400 //-179502.02 * 3.284431e-17 = -5.465239e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010011010011110001011000111101;
		b = 32'b00010110111110010111001000100100;
		correct = 32'b00111011110101001000011100101101;
		#400 //2.6138038e-27 * 4.0300152e-25 = 0.006485841
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101010011111001000111100010011;
		b = 32'b01001110011001101101000010000010;
		correct = 32'b10011011100011000000111011111100;
		#400 //-2.2431735e-13 * 968106100.0 = -2.317074e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010111101110001100011111101101;
		b = 32'b10010010111110100111110100110010;
		correct = 32'b11000100001111001101100010100110;
		#400 //1.194119e-24 * -1.5808081e-27 = -755.38513
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100000100111101101110001011100;
		b = 32'b01010010000001111011100000101010;
		correct = 32'b01001110000101011101001100111110;
		#400 //9.1577e+19 * 145727590000.0 = 628412300.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011001110001000101010110100;
		b = 32'b00001110111100000001000000010110;
		correct = 32'b11111011110001001100101100000111;
		#400 //-12094132.0 * 5.9180058e-30 = -2.0436161e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101100100111111000011010011001;
		b = 32'b01100100111011110000101011001011;
		correct = 32'b11000111001010101101011110111000;
		#400 //-1.5428386e+27 * 3.5276396e+22 = -43735.72
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000101010011101000001101000010;
		b = 32'b10011111101111000101010110100011;
		correct = 32'b01100101000011000101101011001100;
		#400 //-3304.2036 * -7.976277e-20 = 4.142539e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010001010010011111000010010011;
		b = 32'b11100001010110011101001010001111;
		correct = 32'b10101111011011010101010101100000;
		#400 //54207787000.0 * -2.5113224e+20 = -2.1585356e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110110011111001100101010110111;
		b = 32'b01111010011000010110111100111001;
		correct = 32'b00111011100011111000100010001000;
		#400 //1.281807e+33 * 2.9263066e+35 = 0.0043802895
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000001010100111001111000000010;
		b = 32'b00111001101111010100111110010110;
		correct = 32'b01000111000011110001010100000110;
		#400 //13.226076 * 0.00036108185 = 36629.023
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010011110100000001011001001111;
		b = 32'b00010001001100111101110000101100;
		correct = 32'b01000010000101000001011010010110;
		#400 //5.252858e-27 * 1.4188456e-28 = 37.022057
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000010001001010101000010111111;
		b = 32'b01010001101011110010111101011110;
		correct = 32'b00101111111100011001001111010001;
		#400 //41.328854 * 94051746000.0 = 4.3942674e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110100101101011110111011111101;
		b = 32'b11011101110010001101101001110011;
		correct = 32'b11010110011001111110001010110101;
		#400 //1.1531409e+32 * -1.8091258e+18 = -63740220000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101101101100111111001010000001;
		b = 32'b00110010110101010010010011010101;
		correct = 32'b10111010010110000010000011110001;
		#400 //-2.0457637e-11 * 2.4813213e-08 = -0.0008244655
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100110000100001000001011011;
		b = 32'b01110010011100011101111101110111;
		correct = 32'b00010001110011010110011000001010;
		#400 //1552.5111 * 4.7907865e+30 = 3.2406184e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001101111000000101010111110100;
		b = 32'b10101001000000011011001111001101;
		correct = 32'b01100100010111010110010000101111;
		#400 //-470466180.0 * -2.8799706e-14 = 1.6335798e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010100000110110010000110101111;
		b = 32'b00100001100011111010111110010111;
		correct = 32'b01110010000010100011001000111001;
		#400 //2665140200000.0 * 9.736535e-19 = 2.7372574e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000000111110101000010010001010;
		b = 32'b00100101101011011100011001001111;
		correct = 32'b01011010101110001000011100100100;
		#400 //7.828679 * 3.0145095e-16 = 2.5969992e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111101110100110011001110100100;
		b = 32'b11001001011000101100111010101101;
		correct = 32'b00110011111011100110001011000010;
		#400 //-0.10312584 * -929002.8 = 1.11007026e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100111110001101001110101101011;
		b = 32'b00001001001101100001010000101100;
		correct = 32'b11011110000010111001111111110001;
		#400 //-5.5126713e-15 * 2.1916938e-33 = -2.5152563e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010001101001010000110011101011;
		b = 32'b11001100111110110111011011110100;
		correct = 32'b01000100001010000000011011111011;
		#400 //-88610790000.0 * -131839900.0 = 672.1091
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101101001010001100010110010010;
		b = 32'b10101100111000101101110010010001;
		correct = 32'b10111111101111100111001011110100;
		#400 //9.593564e-12 * -6.447794e-12 = -1.4878831
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111001101100101001010010101000;
		b = 32'b10110101010010011111110111110110;
		correct = 32'b01000011111000100101010000111010;
		#400 //-0.00034061563 * -7.5247897e-07 = 452.65802
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110001100100100111110000101110;
		b = 32'b00011111101100011000001011010110;
		correct = 32'b11010001010100110100000101100100;
		#400 //-4.263277e-09 * 7.5178866e-20 = -56708450000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101001010000011001011100110001;
		b = 32'b11010101011100010110110110101111;
		correct = 32'b00010011010011010100011001011101;
		#400 //-4.2985746e-14 * -16590837000000.0 = 2.590933e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010111010100011101110110111001;
		b = 32'b00001101011000110110101001101010;
		correct = 32'b01001001011011000011111010011101;
		#400 //6.7811396e-25 * 7.0077867e-31 = 967657.8
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100110100100011101100011001000;
		b = 32'b11011101011010110010011010111011;
		correct = 32'b00001000100111101100011100010111;
		#400 //-1.0120155e-15 * -1.0590273e+18 = 9.556085e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110100000000100000011111100000;
		b = 32'b10000010100010011101100110011000;
		correct = 32'b01110000111100010111101010100000;
		#400 //-1.2110058e-07 * -2.0255233e-37 = 5.9787306e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000111100011111100111010000;
		b = 32'b10101111110101010010101111111000;
		correct = 32'b01000000100100010100101110101001;
		#400 //-1.7606059e-09 * -3.8775716e-10 = 4.540486
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111100000001001001111011101111;
		b = 32'b10110100010011101110011101101000;
		correct = 32'b11000111001001000001011100100000;
		#400 //0.008094533 * -1.926943e-07 = -42007.125
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011010111111100000011000110101;
		b = 32'b01000001011010101111011011001110;
		correct = 32'b11011001000010100110001000100000;
		#400 //-3.5750734e+16 * 14.685255 = -2434464800000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110100100001010001001101100000;
		b = 32'b01101001100100011000010100001101;
		correct = 32'b01001010011010100001101110111001;
		#400 //8.4346735e+31 * 2.199032e+25 = 3835630.2
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000001111101001111110010000011;
		b = 32'b11111011111110011100100100111011;
		correct = 32'b00000101011110110001010010110111;
		#400 //-30.623297 * -2.5939267e+36 = 1.1805768e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111011101000100101100000110110;
		b = 32'b00001111000000100001011001010010;
		correct = 32'b01101100000111111011110101100110;
		#400 //0.004954363 * 6.4137936e-30 = 7.7245446e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111001101110001010110011000111;
		b = 32'b01011010011011100101000110111111;
		correct = 32'b11011110110001100110000000110010;
		#400 //-1.1986087e+35 * 1.6770231e+16 = -7.14724e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101001010111101110010011101010;
		b = 32'b11101101100001110101101011010001;
		correct = 32'b10111011010100101100100001100111;
		#400 //1.6841409e+25 * -5.2362833e+27 = -0.0032162906
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010010010010010001001000101100;
		b = 32'b00111010100010010011001011101110;
		correct = 32'b01010111001110111001011011101100;
		#400 //215898320000.0 * 0.0010467449 = 206256880000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110100011010100101111100001110;
		b = 32'b11100000101100000110001011110001;
		correct = 32'b00010011001010100001010000010000;
		#400 //-2.1827529e-07 * -1.0167989e+20 = 2.1466908e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110001010110010000000011001111;
		b = 32'b11001010011110000011100111101111;
		correct = 32'b00100110010111111100110010001110;
		#400 //-3.1578116e-09 * -4066939.8 = 7.764589e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011110010001000010110110000101;
		b = 32'b00000101111010010110111110111100;
		correct = 32'b11010111110101110010001111010111;
		#400 //-1.0385567e-20 * 2.195226e-35 = -473097860000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001000010101000101010001000100;
		b = 32'b00001000110101011000000000011100;
		correct = 32'b00111110111111101001100001111000;
		#400 //6.3895483e-34 * 1.284959e-33 = 0.497257
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000001111110000100011001010001;
		b = 32'b11110111101111110110011110101000;
		correct = 32'b10001001101001100000011111110011;
		#400 //31.034334 * -7.7643055e+33 = -3.997052e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000000001011111110000100011001;
		b = 32'b00001011111011101011110001001101;
		correct = 32'b11110011101111001001100100100100;
		#400 //-2.7481139 * 9.195759e-32 = -2.9884579e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011100011101011110100001011101;
		b = 32'b00000110000010111111010100000011;
		correct = 32'b01010101111000001110011000011001;
		#400 //8.1364023e-22 * 2.6323e-35 = 30909858000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000110101110100010001010000001;
		b = 32'b01011001000111101111010110100000;
		correct = 32'b00101101000101011110000111101111;
		#400 //23825.252 * 2796444600000000.0 = 8.519837e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001100011001011011001001000000;
		b = 32'b00100110111111101010100111001000;
		correct = 32'b00100100111001101110011011101011;
		#400 //1.7695158e-31 * 1.767081e-15 = 1.0013779e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001011100100000110010100101011;
		b = 32'b00011000000110101101111100110101;
		correct = 32'b00110010111011101010111010100101;
		#400 //5.5619003e-32 * 2.0016724e-24 = 2.7786266e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001101100001101000100110110111;
		b = 32'b10000100110000000010001100000000;
		correct = 32'b11001000001100110100000110011100;
		#400 //8.291541e-31 * -4.5171125e-36 = -183558.44
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100111111011101101010111110100;
		b = 32'b10000110011100110000100110100110;
		correct = 32'b01100000111110111001001011101111;
		#400 //-6.629024e-15 * -4.571031e-35 = 1.4502251e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010001101010010011000000001100;
		b = 32'b01010101111101010011001001001010;
		correct = 32'b10111011001100001010010001101001;
		#400 //-90831946000.0 * 33699542000000.0 = -0.0026953465
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111111111010011010011000111100;
		b = 32'b11110001101100000100011001100001;
		correct = 32'b10001101101010011010100101101011;
		#400 //1.8253856 * -1.7457422e+30 = -1.0456215e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010101101010111101011111110100;
		b = 32'b00111101110011011011111001011110;
		correct = 32'b01010111010101011101000110111100;
		#400 //23618000000000.0 * 0.10046075 = 235096780000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011100110010100111100111000001;
		b = 32'b01101001001101000110110111000111;
		correct = 32'b10110011000011111010001111110101;
		#400 //-4.5593452e+17 * 1.3632816e+25 = -3.34439e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111001101111000011001100011000;
		b = 32'b10100101111101011101011000001000;
		correct = 32'b01010011010000111111101100000111;
		#400 //-0.00035896222 * -4.2645758e-16 = 841730160000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011011110100011010101001110011;
		b = 32'b10101011111101011011011010010100;
		correct = 32'b11101111010110100111000110001001;
		#400 //1.1803136e+17 * -1.7458973e-12 = -6.760499e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010000100111010100111110000011;
		b = 32'b01001011001100001100111011110111;
		correct = 32'b00000100111000111100010011100111;
		#400 //6.204809e-29 * 11587319.0 = 5.354827e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101010010011000011000011101111;
		b = 32'b11010000110011000011011010010100;
		correct = 32'b01011000111111111111100011101101;
		#400 //-6.1712987e+25 * -27409031000.0 = 2251556700000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010011010011011111010110010011;
		b = 32'b00001010111101100110001000000011;
		correct = 32'b11000111110101011111111110100001;
		#400 //-2.5995715e-27 * 2.3725806e-32 = -109567.26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010011010011011001100001110010;
		b = 32'b00100010111011010001111110111010;
		correct = 32'b00101111110111011111011000110110;
		#400 //2.5949799e-27 * 6.427257e-18 = 4.037461e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001001100001000001100110001011;
		b = 32'b01111011100110000101010110001011;
		correct = 32'b00001101010111011111111011101101;
		#400 //1082161.4 * 1.5819283e+36 = 6.840774e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101110100111100010001100000111;
		b = 32'b11100100110101101101100000011001;
		correct = 32'b00001001001111000110111000000101;
		#400 //-7.19123e-11 * -3.1705398e+22 = 2.2681408e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011001100100101010100101110100;
		b = 32'b00100111100001010101100011110001;
		correct = 32'b11110001100011001100011111010011;
		#400 //-5160208000000000.0 * 3.7011346e-15 = -1.3942232e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001010101001001011101111110011;
		b = 32'b00011001101111010011001010100110;
		correct = 32'b10110000010111101110011000010000;
		#400 //-1.5863324e-32 * 1.9562599e-23 = -8.109007e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100111100000110001011110110010;
		b = 32'b11100101101001010100101100110111;
		correct = 32'b01000001010010110000011111010011;
		#400 //-1.2381342e+24 * -9.757224e+22 = 12.68941
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000111111100000001010011010010;
		b = 32'b00111010100111010000101001001001;
		correct = 32'b11001100110000111010111101011110;
		#400 //-122921.64 * 0.0011981215 = -102595310.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101101001010100001011000011000;
		b = 32'b10111101100110001010010010000001;
		correct = 32'b00101111000011101010000010101010;
		#400 //-9.668287e-12 * -0.07453252 = 1.2971904e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111011101101000011110111101011;
		b = 32'b10110101101101010000100011110101;
		correct = 32'b11000101011111101110000011100010;
		#400 //0.0055005453 * -1.3488158e-06 = -4078.0552
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101010110010101110101011011110;
		b = 32'b01001001111111001101111001110010;
		correct = 32'b01100000010011010110111000010101;
		#400 //1.2265607e+26 * 2071502.2 = 5.921117e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110010001101010101101111001000;
		b = 32'b01110011111111000110100110110001;
		correct = 32'b00111101101101111110111110010110;
		#400 //3.5921756e+30 * 3.9996414e+31 = 0.08981244
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000100000111001110101001110100;
		b = 32'b01110000101000111100101100100111;
		correct = 32'b10010010111101010100000000100001;
		#400 //-627.6633 * 4.0553322e+29 = -1.5477483e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100011111011010010000011011000;
		b = 32'b10110101011010101010110111100000;
		correct = 32'b01101110000000010101010111110111;
		#400 //-8.74849e+21 * -8.7424814e-07 = 1.0006873e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101100001000000010001111011010;
		b = 32'b01100111100011100001100010101101;
		correct = 32'b10000100000100000100000011110001;
		#400 //-2.275727e-12 * 1.3420625e+24 = -1.6956938e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110010100101110101100011110011;
		b = 32'b10001111111011100100011011010110;
		correct = 32'b11100010001000101001101011011000;
		#400 //1.7619163e-08 * -2.3495897e-29 = -7.4988255e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101011011001001010010010101010;
		b = 32'b11010010110010000001100101000110;
		correct = 32'b01011000000100100100001001101100;
		#400 //-2.764127e+26 * -429708740000.0 = 643255900000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001000100101000011001011110111;
		b = 32'b00101101000000001100000011110010;
		correct = 32'b11011011000100110101010011100001;
		#400 //-303511.72 * 7.3188e-12 = -4.1470147e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110111110010100101010011100000;
		b = 32'b10110000001110101100001100110011;
		correct = 32'b11000111000010101010101110100010;
		#400 //2.41198e-05 * -6.79438e-10 = -35499.633
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101101000000001101000011010011;
		b = 32'b11101000001101101000000100001001;
		correct = 32'b11000100001101001011000011100000;
		#400 //2.4916584e+27 * -3.447404e+24 = -722.7637
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010101111010000110110000010000;
		b = 32'b00101010000100000000101001011101;
		correct = 32'b01101011010011101000101000010101;
		#400 //31943853000000.0 * 1.2793365e-13 = 2.496908e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111100001011000010110110101011;
		b = 32'b11110111110111011110111100100111;
		correct = 32'b01000011110001101001101101100000;
		#400 //-3.5760053e+36 * -9.00272e+33 = 397.21387
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001000111001000011100011101000;
		b = 32'b01111000101111001001111001010100;
		correct = 32'b10001111100110101110000000111010;
		#400 //-467399.25 * 3.0605096e+34 = -1.5271941e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011110001010110011011000010011;
		b = 32'b01011001011000000010111011011010;
		correct = 32'b01000100010000111000001010011111;
		#400 //3.0842673e+18 * 3943869300000000.0 = 782.04095
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101001100011001100101010111111;
		b = 32'b01110010101111111100101000110010;
		correct = 32'b00110110001110111110110110101001;
		#400 //2.1275882e+25 * 7.597578e+30 = 2.8003508e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111110011111101000001101011111;
		b = 32'b11100011001001011000000000101100;
		correct = 32'b01011010110001001101011111011101;
		#400 //-8.4576507e+37 * -3.0529485e+21 = 2.770322e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001101100001010101001000001000;
		b = 32'b10011000011111000000000000011010;
		correct = 32'b00110100100001110110111110111001;
		#400 //-8.216506e-31 * -3.2570288e-24 = 2.5226998e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110011111111000001011111110101;
		b = 32'b00111010000101110011111100110010;
		correct = 32'b10111001010101010101100010110000;
		#400 //-1.1739022e-07 * 0.00057696097 = -0.00020346302
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000000010101101000011001001110;
		b = 32'b00001001101010011110010101111010;
		correct = 32'b00110110000000100110000000011000;
		#400 //7.946032e-39 * 4.090107e-33 = 1.9427443e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111111011000000011000110100111;
		b = 32'b11010101011010010010100110000001;
		correct = 32'b11101001011101100010011101000110;
		#400 //2.9800488e+38 * -16022779000000.0 = -1.8598826e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010110111010111010111111110111;
		b = 32'b00100001110001110100000110000001;
		correct = 32'b11110100100101110110011100111010;
		#400 //-129570500000000.0 * 1.3502103e-18 = -9.59632e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001000101011110100001101111000;
		b = 32'b10111010010110010011001101001101;
		correct = 32'b00001101110011101001001001011111;
		#400 //-1.0548291e-33 * -0.00082855375 = 1.2730968e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000000010110110101111000100001;
		b = 32'b10101111011010010010001111011010;
		correct = 32'b01010000011100001110000010010010;
		#400 //-3.4276202 * -2.1203964e-10 = 16164997000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000111011101011011100111001110;
		b = 32'b10111001010010111110000100010101;
		correct = 32'b01001101100110100100010110110001;
		#400 //-62905.805 * -0.00019443438 = 323532320.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000101111111111111010001011110;
		b = 32'b01101110011101000011010001000010;
		correct = 32'b00010111000001100010100010110101;
		#400 //8190.546 * 1.889438e+28 = 4.3349115e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011000101001101011100001010110;
		b = 32'b01001011101010011111110010111001;
		correct = 32'b10001100011110110001010001101000;
		#400 //-4.3096126e-24 * 22280562.0 = -1.9342477e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011011011101011010101011110001;
		b = 32'b01011010001011000110000001110010;
		correct = 32'b01000000101101100110110001000101;
		#400 //6.914932e+16 * 1.2129935e+16 = 5.7007165
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010010010010000010001001000000;
		b = 32'b10111001011011101100100000101000;
		correct = 32'b01011000010101101001000010101001;
		#400 //-214892020000.0 * -0.00022772013 = 943667200000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111001011011111001001111000110;
		b = 32'b00001110010110010110001100111010;
		correct = 32'b01101010100011010001000011000011;
		#400 //0.00022847866 * 2.679509e-30 = 8.526885e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001001110011010011111011111111;
		b = 32'b00101000011001101100101101111011;
		correct = 32'b11100000111000111010100100111010;
		#400 //-1681375.9 * 1.28116876e-14 = -1.31237655e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101111011011011000001011111000;
		b = 32'b11011010111110010100001111100111;
		correct = 32'b11010011111100111110110111000101;
		#400 //7.350628e+28 * -3.5080964e+16 = -2095332300000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101100001010110010101000011111;
		b = 32'b00111000110001111111111011011101;
		correct = 32'b10110010110110110001100001110001;
		#400 //-2.4323943e-12 * 9.5365314e-05 = -2.550607e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010001110100011111101111100001;
		b = 32'b10111110111000010010000010010000;
		correct = 32'b10010010011011101100011110110000;
		#400 //3.3129618e-28 * -0.43970156 = -7.534569e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011000010001101011111011000100;
		b = 32'b01001101101110010000001100000110;
		correct = 32'b10001010000010011000000001011100;
		#400 //-2.5687212e-24 * 387997900.0 = -6.620452e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000110101011101110001000100100;
		b = 32'b00101101000001101010100111011100;
		correct = 32'b00011001001001100011101011001011;
		#400 //6.578381e-35 * 7.6547345e-12 = 8.593872e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101111100100110001101000110111;
		b = 32'b11011111111001000111101001010101;
		correct = 32'b01001111001001001101001001111001;
		#400 //-9.105198e+28 * -3.292713e+19 = 2765257000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100100110001011100110101100000;
		b = 32'b01011011010001111101110100101101;
		correct = 32'b00001000111111010101101111110101;
		#400 //8.578305e-17 * 5.6256706e+16 = 1.5248503e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001010101100011001000001101101;
		b = 32'b00011111111000011110011110101000;
		correct = 32'b11101010010010010011100000100100;
		#400 //-5818422.5 * 9.567445e-20 = -6.08148e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010111001110000001001111100010;
		b = 32'b00000011101100000000011110001110;
		correct = 32'b11010011000001011101101000101011;
		#400 //-5.94787e-25 * 1.0346085e-36 = -574890900000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000101001111101001001111111100;
		b = 32'b11011011001000111010100101000010;
		correct = 32'b00101001100101010000110101000011;
		#400 //-3049.249 * -4.606652e+16 = 6.61923e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011101010111000010101111000101;
		b = 32'b11010101001000000111000101101110;
		correct = 32'b01000111101011111010011001111110;
		#400 //-9.915619e+17 * -11025565000000.0 = 89932.984
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111111011100101000110011010011;
		b = 32'b01101001000111010111110100010111;
		correct = 32'b11010101110001010010001001100010;
		#400 //-3.2240438e+38 * 1.1899505e+25 = -27093933000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101010011010001110110011010101;
		b = 32'b11110100011101000001011011011110;
		correct = 32'b00110101011101000100101010000001;
		#400 //-7.03973e+25 * -7.7354995e+31 = 9.10055e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101110001010110011000000100101;
		b = 32'b10100010101011100100010011111010;
		correct = 32'b11001010111110110111100100110111;
		#400 //3.892366e-11 * -4.7235826e-18 = -8240283.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001101110011011101111110100111;
		b = 32'b00101010011010011110011000111111;
		correct = 32'b10100010111000010101001101111111;
		#400 //-1.2687943e-30 * 2.077444e-13 = -6.1074777e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110010011110001010101011110011;
		b = 32'b11011101110000010010111001000001;
		correct = 32'b00010100001001001100001111101011;
		#400 //-1.4474369e-08 * -1.7400169e+18 = 8.318522e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001010010110001100101101100101;
		b = 32'b10001010010111000000111101010101;
		correct = 32'b00111111011111000011001110001010;
		#400 //-1.0438276e-32 * -1.0595498e-32 = 0.9851614
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100110101111110100110011110001;
		b = 32'b11100100111000111010010000011100;
		correct = 32'b11000001010101110010000111011110;
		#400 //4.5169566e+23 * -3.359389e+22 = -13.445768
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010100001111011101111011100011;
		b = 32'b10111101000100001110001100101110;
		correct = 32'b10010110101001111011110101111101;
		#400 //9.586018e-27 * -0.035372905 = -2.709989e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001001011111001001010100100001;
		b = 32'b11001001100001010010000001010000;
		correct = 32'b00111111011100101101101101000010;
		#400 //-1034578.06 * -1090570.0 = 0.9486581
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000000011000001000000110100000;
		b = 32'b00110110001110010001111110010111;
		correct = 32'b01001001100110110011101100000111;
		#400 //3.5079117 * 2.7585536e-06 = 1271648.9
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110100111111111010111001110100;
		b = 32'b01000011110011011001100101100100;
		correct = 32'b10110000100111110010111000000100;
		#400 //-4.7624383e-07 * 411.19836 = -1.1581851e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100010011000011000010000000011;
		b = 32'b00100011010000101000011011011001;
		correct = 32'b11111110100101000110010000010100;
		#400 //-1.0400075e+21 * 1.0545316e-17 = -9.862269e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000110111010110100000100010000;
		b = 32'b00110110010010111100001111111001;
		correct = 32'b00010000000100111100011111000010;
		#400 //8.8492776e-35 * 3.0363428e-06 = 2.9144526e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001100111111110010110000110110;
		b = 32'b11001011111111101100101010101100;
		correct = 32'b00000000100000000011000100000000;
		#400 //-3.931558e-31 * -33396056.0 = 1.1772521e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100110011111011000000100110100;
		b = 32'b01100000111011100011000111101110;
		correct = 32'b11000101000010000011101000011110;
		#400 //-2.9928552e+23 * 1.3731009e+20 = -2179.6323
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100110010000010000011000011010;
		b = 32'b00110010001100001011000101111111;
		correct = 32'b10110011100010111101010010000010;
		#400 //-6.6968595e-16 * 1.0284906e-08 = -6.511347e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100110110110100001110010001001;
		b = 32'b11011000001110110100000100100010;
		correct = 32'b01001110000101010001011110111011;
		#400 //-5.1500114e+23 * -823553700000000.0 = 625340100.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111011000000011100100111111011;
		b = 32'b10110000101010101000011001001110;
		correct = 32'b01001001110000101101100001111100;
		#400 //-0.0019804228 * -1.24073e-09 = 1596175.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101101010110011111011011011101;
		b = 32'b01100110100001111010100000010010;
		correct = 32'b11000110010011011010100110001100;
		#400 //-4.216043e+27 * 3.203099e+23 = -13162.387
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011011100100110111100101001000;
		b = 32'b01100011010011000001111110000011;
		correct = 32'b10110111101110001111010000011001;
		#400 //-8.302034e+16 * 3.7654064e+21 = -2.2048176e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011100111000101100011001110100;
		b = 32'b10011001000100110011001011010010;
		correct = 32'b01000011010001010011001010100100;
		#400 //-1.5006724e-21 * -7.609985e-24 = 197.19781
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011011000111001011011110010111;
		b = 32'b10011011001111000010101110100011;
		correct = 32'b10111111010101010011010101110001;
		#400 //1.2963339e-22 * -1.5565095e-22 = -0.8328467
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111000000010100101001000101111;
		b = 32'b00101010001010100101100111010000;
		correct = 32'b11001101010011111101110111000001;
		#400 //-3.2978303e-05 * 1.5130193e-13 = -217963540.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111001100110010100001010010100;
		b = 32'b01100111000010101110000010110010;
		correct = 32'b00010010000011010100000101111111;
		#400 //0.0002923204 * 6.558315e+23 = 4.4572485e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111111010101010011110110100100;
		b = 32'b01111101000101011100100101101100;
		correct = 32'b11000001101101100011100101110111;
		#400 //-2.8344562e+38 * 1.2443801e+37 = -22.778059
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100110001111101100011011111100;
		b = 32'b11000000010111101110101000100101;
		correct = 32'b00100101010110110001011111000000;
		#400 //-6.6189166e-16 * -3.483041 = 1.9003269e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100100000001010011001010100111;
		b = 32'b11011001111010010001101101001110;
		correct = 32'b00001001100100100100011101111001;
		#400 //-2.8882682e-17 * -8201711400000000.0 = 3.5215434e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100010111011100001011110101111;
		b = 32'b00000011001110110001100000110011;
		correct = 32'b11011111001000101110001111011100;
		#400 //-6.4535105e-18 * 5.498214e-37 = -1.1737467e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101100111001100110010110101101;
		b = 32'b11010101110101010000010100000001;
		correct = 32'b00010110100010100111000100100011;
		#400 //-6.5482814e-12 * -29277184000000.0 = 2.2366502e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000001101011111001001110101010;
		b = 32'b11001100110100111011010000011100;
		correct = 32'b00110100010101000101000001101101;
		#400 //-21.947102 * -110993630.0 = 1.9773297e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110110001100000001111011111011;
		b = 32'b11010101010001100001001010010101;
		correct = 32'b01100000011000111010000011101010;
		#400 //-8.9303965e+32 * -13611444000000.0 = 6.560947e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101001110011110001011001111000;
		b = 32'b00111011100001111111011101000100;
		correct = 32'b00101101110000101111010001111110;
		#400 //9.1965444e-14 * 0.0041493494 = 2.2163823e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101101011010110110100111010011;
		b = 32'b00011110101010111101100001010110;
		correct = 32'b01001110001011110101100101101100;
		#400 //1.3381701e-11 * 1.8194804e-20 = 735468300.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011011011111000110000010010111;
		b = 32'b00011110011111100110100111111111;
		correct = 32'b11111100011111011111001101011000;
		#400 //-7.1037896e+16 * 1.34685675e-20 = -5.2743468e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000110100110111011001001100010;
		b = 32'b11011101111011110001000011011000;
		correct = 32'b10101000001001101011100110111111;
		#400 //19929.191 * -2.1533133e+18 = -9.255128e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011110001010000100101001010110;
		b = 32'b00111011110110110011110101100111;
		correct = 32'b01100001110001001000000111111110;
		#400 //3.03165e+18 * 0.0066906693 = 4.531161e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001100101100011100000110011001;
		b = 32'b01001011110010011000110010011111;
		correct = 32'b11000000011000011100011101101100;
		#400 //-93195464.0 * 26417470.0 = -3.5277967
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110110101000100001001100000010;
		b = 32'b00111000101110010111001110010011;
		correct = 32'b11111101010111111011101011010000;
		#400 //-1.6436282e+33 * 8.843015e-05 = -1.8586739e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001010101111011100110101000001;
		b = 32'b00010100000101010001000000100000;
		correct = 32'b10110110001000101111101101110111;
		#400 //-1.8277246e-32 * 7.525758e-27 = -2.4286253e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011010101000100110100111011111;
		b = 32'b00110101011001011110110111100110;
		correct = 32'b00100100101101001101010000110110;
		#400 //6.7172674e-23 * 8.5655336e-07 = 7.8422056e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001001110001111110101010101011;
		b = 32'b10011000101000101110100110011111;
		correct = 32'b10110000100111010001001011110011;
		#400 //4.8128188e-33 * -4.2111916e-24 = -1.1428639e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011101100111110000101010110011;
		b = 32'b10101110011101110111100010101000;
		correct = 32'b11101110101001001000010111011101;
		#400 //1.4325211e+18 * -5.6268462e-11 = -2.5458686e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010001101100110101100000000011;
		b = 32'b00010011000001101111010101100110;
		correct = 32'b00111110001010100001100010111111;
		#400 //2.8295462e-28 * 1.7034169e-27 = 0.16611002
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111101111110010110110111001101;
		b = 32'b11111100100111011110001100110010;
		correct = 32'b01000000110010100011011010000111;
		#400 //-4.1443486e+37 * -6.5583894e+36 = 6.319156
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111001100111011010101100001011;
		b = 32'b01110000010000111110111101110000;
		correct = 32'b11001000110011100000000001111100;
		#400 //-1.0233247e+35 * 2.4255616e+29 = -421891.88
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001011100100010101110000111010;
		b = 32'b10111010100110000001001011111110;
		correct = 32'b00010000011101001011001010100110;
		#400 //-5.5990735e-32 * -0.001160234 = 4.825814e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110000111000100100010011001010;
		b = 32'b11111010100010101000010000100101;
		correct = 32'b10110101110100010001011100011111;
		#400 //5.602142e+29 * -3.596086e+35 = -1.5578443e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111010010100011010101111100011;
		b = 32'b11110000001111000010101010100010;
		correct = 32'b01001001100011101010000011110001;
		#400 //-2.7216908e+35 * -2.3293889e+29 = 1168414.1
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110100100110111110100010010010;
		b = 32'b10101101111001001110010010010100;
		correct = 32'b11000110001011100101111101001101;
		#400 //2.9040217e-07 * -2.6022108e-11 = -11159.825
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111111111000011100100010101010;
		b = 32'b00011111011100000001010001111010;
		correct = 32'b11011111111100001100000110000000;
		#400 //-1.7639363 * 5.0838915e-20 = -3.4696576e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101001111101110100101010101001;
		b = 32'b11001011000000110011010111001110;
		correct = 32'b00011110011100010011110111001110;
		#400 //-1.0981955e-13 * -8598990.0 = 1.2771215e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011111010001100011101001101101;
		b = 32'b00001111101101110010110111110011;
		correct = 32'b11001111000010101000001111111101;
		#400 //-4.197646e-20 * 1.8062892e-29 = -2323905800.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001011101110000001000010000110;
		b = 32'b10101000110101110101010011000111;
		correct = 32'b11100010010110101101010000000011;
		#400 //24125708.0 * -2.3906561e-14 = -1.0091668e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111110011010010110101000010110;
		b = 32'b11011011101001100000110011011000;
		correct = 32'b00100010001100111110110110000101;
		#400 //-0.22794375 * -9.347794e+16 = 2.4384765e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001010100111011101100010010001;
		b = 32'b00110101001110110100100001110010;
		correct = 32'b11010100110101111100001100010111;
		#400 //-5172296.5 * 6.976835e-07 = -7413528300000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110111010110101010001111111010;
		b = 32'b11000001101001111010110000110010;
		correct = 32'b11110101001001101110100010010011;
		#400 //4.434557e+33 * -20.95908 = -2.1158165e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000110001001001111001111111101;
		b = 32'b10101010111011000100100011001100;
		correct = 32'b10011010101100101011011110000001;
		#400 //3.1024226e-35 * -4.1972534e-13 = -7.391554e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001010011111110101011011011000;
		b = 32'b11000101101110001010001000100110;
		correct = 32'b00000100001100010000010010010111;
		#400 //-1.2294137e-32 * -5908.2686 = 2.0808358e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010000111111001001011101010111;
		b = 32'b00111010111110000110100110000100;
		correct = 32'b01010101100000100010011101000000;
		#400 //33902213000.0 * 0.0018952345 = 17888136000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011111110000001001010111111000;
		b = 32'b11001101111101100011100001100000;
		correct = 32'b01010001010010000011110000111010;
		#400 //-2.775454e+19 * -516361200.0 = 53750243000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111110110011001111111101001101;
		b = 32'b00110010110101110011111001111111;
		correct = 32'b11001011011100111101000000011100;
		#400 //-0.4003853 * 2.5057714e-08 = -15978524.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110100011101100110111111111110;
		b = 32'b10011010001101111100101111111100;
		correct = 32'b11011001101010111001111111010001;
		#400 //2.2951278e-07 * -3.800829e-23 = -6038492600000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011010001111111111111011101100;
		b = 32'b01011100011101110000111001111010;
		correct = 32'b00111101010001101111001000110000;
		#400 //1.3510503e+16 * 2.7816095e+17 = 0.04857081
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101010010101011010100101000101;
		b = 32'b00010110000011110010011001101000;
		correct = 32'b11010011101111110000110001111100;
		#400 //-1.8976928e-13 * 1.1563567e-25 = -1641096400000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001000111011100110001111101111;
		b = 32'b10001111010111111001011000110111;
		correct = 32'b01111001000010000111100110001110;
		#400 //-488223.47 * -1.1023679e-29 = 4.428861e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100001010111001010010000001010;
		b = 32'b11000100000110011010100001110100;
		correct = 32'b11011100101101111100110001000010;
		#400 //2.543815e+20 * -614.6321 = -4.1387604e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000000010101110001001100010110;
		b = 32'b01011000111111101110101110011111;
		correct = 32'b00100110110101111111110001000100;
		#400 //3.36054 * 2242303500000000.0 = 1.4986999e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001110001010100100001110111001;
		b = 32'b00111010111110010110011110000001;
		correct = 32'b01010010101011101100010001101111;
		#400 //714141250.0 * 0.0019028039 = 375309960000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011100011110010100101101101111;
		b = 32'b11011110100101010000100110111101;
		correct = 32'b00111101010101100001101011000001;
		#400 //-2.8068084e+17 * -5.3696613e+18 = 0.05227161
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110101111001111011101001001;
		b = 32'b01101111001011000111000110011110;
		correct = 32'b10000111000011000100001110001111;
		#400 //-5.6316244e-06 * 5.3368776e+28 = -1.0552283e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101100011100011001010010000101;
		b = 32'b10001110001110011011100001000010;
		correct = 32'b11011101101001100111111111100100;
		#400 //3.4330605e-12 * -2.2891727e-30 = -1.4996948e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000001000011110111101110111111;
		b = 32'b00110010010000000010001110011001;
		correct = 32'b11001110001111110010110000111000;
		#400 //-8.967711 * 1.1183965e-08 = -801836540.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100001101100100011010110111011;
		b = 32'b00100001110011110010001101010101;
		correct = 32'b10111111010111000011111101111100;
		#400 //-1.2075972e-18 * 1.4036218e-18 = -0.8603437
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000000101111101001011110001100;
		b = 32'b10001100101110101101010000111010;
		correct = 32'b10110011100000101001001111111101;
		#400 //1.7503109e-38 * -2.8785567e-31 = -6.080516e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000101011110101011000110101001;
		b = 32'b00101011000001101001001101000001;
		correct = 32'b11011001111011100111001000000001;
		#400 //-4011.1038 * 4.781072e-13 = -8389549000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000000101001011000011110001000;
		b = 32'b00111011000011101011000100111100;
		correct = 32'b00000101000101000111110001010101;
		#400 //1.5201476e-38 * 0.002177312 = 6.981763e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010111101010110010111101000001;
		b = 32'b10010100111100100100111001001000;
		correct = 32'b11000010001101001101101111111011;
		#400 //1.1062545e-24 * -2.4466632e-26 = -45.214825
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101001010001000101110101111000;
		b = 32'b01001010111000110000010111100001;
		correct = 32'b10011101110111010110110111010011;
		#400 //-4.3601814e-14 * 7439088.5 = -5.861177e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101111110110011110111000100000;
		b = 32'b01011110001001000011010100110010;
		correct = 32'b00010001001010011110000001101001;
		#400 //3.9641268e-10 * 2.9581046e+18 = 1.3400901e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110010110011001011011110111101;
		b = 32'b10000011111100000010111111100100;
		correct = 32'b11101110010110100011001000001100;
		#400 //2.383228e-08 * -1.4116927e-36 = -1.6882059e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100101111110011110001010101110;
		b = 32'b11010101000101101001011010111101;
		correct = 32'b11010000010101000110011011011110;
		#400 //1.47506345e+23 * -10348385000000.0 = -14254045000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110101110001110111001101010110;
		b = 32'b10111001111110100011111100001001;
		correct = 32'b01111011010011000000100101010000;
		#400 //-5.0566717e+32 * -0.0004773068 = 1.0594174e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101101111011001101011001010010;
		b = 32'b11110001111110101011111101000001;
		correct = 32'b00111011011100011100110001111000;
		#400 //-9.162195e+27 * -2.4832789e+30 = 0.0036895555
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000010111010011101110001001101;
		b = 32'b01100001110011110000001001011111;
		correct = 32'b10100000100100001001101001011011;
		#400 //-116.930275 * 4.7733086e+20 = -2.4496693e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011101110010111100100110001000;
		b = 32'b01101111000000001000111110000011;
		correct = 32'b10101110010010101110011000001011;
		#400 //-1.8355522e+18 * 3.9787576e+28 = -4.61338e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111001001011000010000110100100;
		b = 32'b00011110100110111010000111000011;
		correct = 32'b11011010000011011001000111110010;
		#400 //-0.0001641573 * 1.6478166e-20 = -9962110000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011000111111111000010011000000;
		b = 32'b00101011000101110001110000001001;
		correct = 32'b10101101010110000111000100001001;
		#400 //-6.605e-24 * 5.3684883e-13 = -1.2303277e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110010001110001000001011101111;
		b = 32'b10001010001110101010101011010111;
		correct = 32'b11100111011111010000101100011010;
		#400 //1.07399805e-08 * -8.987706e-33 = -1.1949635e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010100111101101001001110111011;
		b = 32'b10101010000100000100001010111111;
		correct = 32'b11101010010110101100100010010011;
		#400 //8472323700000.0 * -1.2812926e-13 = -6.6123253e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001100100001100010010111111101;
		b = 32'b10100100010111100011010101110110;
		correct = 32'b10100111100110101000110001011011;
		#400 //2.0668832e-31 * -4.818386e-17 = -4.289576e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101101100101111110111100001100;
		b = 32'b10011101010101100101010111000100;
		correct = 32'b11001111101101010111011111101101;
		#400 //1.727287e-11 * -2.8367004e-21 = -6089071000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000100100101010110100100001111;
		b = 32'b01011000110001100101101000011100;
		correct = 32'b10101011010000001101010110010010;
		#400 //-1195.2831 * 1744722600000000.0 = -6.850849e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010110000111000111110101110;
		b = 32'b10110010100111111011000100100111;
		correct = 32'b01000111100111001100000000110001;
		#400 //-0.0014920139 * -1.8590596e-08 = 80256.38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100100101101011110100101100011;
		b = 32'b01000111101111000100110010101111;
		correct = 32'b11011100011101110101000011000001;
		#400 //-2.6845424e+22 * 96409.37 = -2.7845244e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011010011000100111111001010001;
		b = 32'b11010110010101000000100000010011;
		correct = 32'b11000011100010001011101011111100;
		#400 //1.5938058e+16 * -58282786000000.0 = -273.46082
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011110000011010011011101111101;
		b = 32'b01110100000110001001100111011000;
		correct = 32'b00101001011011001110011011110001;
		#400 //2.5439348e+18 * 4.836117e+31 = 5.2602837e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001010100101111111011101110010;
		b = 32'b11100010110100010101101010100000;
		correct = 32'b10100111001110011101001101111110;
		#400 //4979641.0 * -1.9309499e+21 = -2.5788558e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101101001000110101001011100111;
		b = 32'b11111011011100010111000001011001;
		correct = 32'b10110001001011010010110010000011;
		#400 //3.1591425e+27 * -1.2536222e+36 = -2.5200115e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100000011011011010111110001001;
		b = 32'b00001100111100110001001000010111;
		correct = 32'b11010010111110100101010000011110;
		#400 //-2.013276e-19 * 3.7450966e-31 = -537576540000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111001000000101100101110110000;
		b = 32'b01101010000000101011111110001001;
		correct = 32'b11001110100000000000101111100110;
		#400 //-4.2445617e+34 * 3.9516214e+25 = -1074131700.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111010101010100111011001011101;
		b = 32'b11010111010010101100010011101111;
		correct = 32'b11100010110101110011011001000000;
		#400 //4.4254558e+35 * -222947170000000.0 = -1.9849796e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010000011111011100110110011011;
		b = 32'b11011011011100101111100101011010;
		correct = 32'b00110100100001011011010001110000;
		#400 //-17032441000.0 * -6.839111e+16 = 2.4904466e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110111101010000111111110000101;
		b = 32'b10001100010011101101001111111000;
		correct = 32'b11101010110100001000111010110101;
		#400 //2.0086542e-05 * -1.593345e-31 = -1.2606524e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101111001000011111110010010111;
		b = 32'b11101100111011111111101001110110;
		correct = 32'b10000001101011001100110100100111;
		#400 //1.4732603e-10 * -2.3209283e+27 = -6.34772e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111000000011110000110011000010;
		b = 32'b11011101100000101101111011100100;
		correct = 32'b11011010000010111110100101111010;
		#400 //1.1605581e+34 * -1.1787782e+18 = -9845433000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000110111100010111010100000001;
		b = 32'b00010101111111101111101000010100;
		correct = 32'b01110000011100100110110100001010;
		#400 //30906.502 * 1.02984337e-25 = 3.0010877e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011000100000011000101111001111;
		b = 32'b01000011011000100110000001010111;
		correct = 32'b10010100100100100111111110100010;
		#400 //-3.348689e-24 * 226.37633 = -1.4792575e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011111100110001101101010011110;
		b = 32'b10010001110111110011111000000000;
		correct = 32'b01001101001011110100100010000011;
		#400 //-6.4736176e-20 * -3.5221407e-28 = 183797810.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100111010001000010101001100110;
		b = 32'b10101001011110001110110111111111;
		correct = 32'b01111101010010011011110010111111;
		#400 //-9.2636594e+23 * -5.527349e-14 = 1.6759678e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011111111000010001010110000011;
		b = 32'b01010101101001001010011111001101;
		correct = 32'b00001001101011101111100111011011;
		#400 //9.5326795e-20 * 22630076000000.0 = 4.212394e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111001010110000010001101111000;
		b = 32'b10010001000110100001011001101001;
		correct = 32'b01100111101100111000101110101010;
		#400 //-0.00020612578 * -1.2155364e-28 = 1.6957599e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001000111100011110100011100100;
		b = 32'b11001000000110001010101000100010;
		correct = 32'b11000000010010101101001110011111;
		#400 //495431.12 * -156328.53 = -3.1691663
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110101001011100111111101110100;
		b = 32'b10111010101010010100001111010010;
		correct = 32'b11111010000000111111010100001100;
		#400 //2.2120232e+32 * -0.0012913889 = -1.7129026e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110011110110011101100110000001;
		b = 32'b00100100011001000110111000011101;
		correct = 32'b01001110111101000010010001111011;
		#400 //1.0144414e-07 * 4.953289e-17 = 2048015700.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011000010110000100011100111000;
		b = 32'b00011111010111110110010001010010;
		correct = 32'b00111000011101111101100100010011;
		#400 //2.7953302e-24 * 4.730507e-20 = 5.9091555e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000110011010010001101101111010;
		b = 32'b01100101000100111000101110010101;
		correct = 32'b00100000110010100011101001001100;
		#400 //14918.869 * 4.354767e+22 = 3.4258709e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110010111111100111101110011100;
		b = 32'b00000010111100010001001110001010;
		correct = 32'b11101111100001110001111001000100;
		#400 //-2.9625703e-08 * 3.5422982e-37 = -8.363413e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100001011001111100010001001000;
		b = 32'b10010110111010000000101001110111;
		correct = 32'b11001001111111111011001010010010;
		#400 //7.852562e-19 * -3.7488226e-25 = -2094674.2
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110010100001111001101111100;
		b = 32'b11110101111001001100010001001101;
		correct = 32'b10000111111010011101001101001100;
		#400 //0.20405382 * -5.7999274e+32 = -3.5182133e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010110010111001100101110011101;
		b = 32'b10111101010101111100011001101000;
		correct = 32'b10011000100000101111101001100110;
		#400 //1.7835707e-25 * -0.05267945 = -3.385705e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010010111111011100000010011111;
		b = 32'b11100011100011000111101011110100;
		correct = 32'b10101110111001110011010110000011;
		#400 //544929200000.0 * -5.182808e+21 = -1.05141694e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100111011100000010000101000101;
		b = 32'b00011001111111100011000001001111;
		correct = 32'b01001100111100011101011101010001;
		#400 //3.3324726e-15 * 2.6282496e-23 = 126794376.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111011111011110101100000001101;
		b = 32'b11010010010011111011100010100011;
		correct = 32'b11101001000100110111110001111011;
		#400 //2.4854897e+36 * -223038980000.0 = -1.1143746e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001110011100001100001011010011;
		b = 32'b10100011001110110000100001011010;
		correct = 32'b11101010101001001100010100101111;
		#400 //1009824960.0 * -1.0139059e-17 = -9.95975e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100100000111000001001010110000;
		b = 32'b10000100000110000000001101000100;
		correct = 32'b11011111100000110110101100111011;
		#400 //3.3842937e-17 * -1.7869014e-36 = -1.8939455e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100001000000110001111010001010;
		b = 32'b00001101100011101110010111001001;
		correct = 32'b11010010111010101110011000110101;
		#400 //-4.4424945e-19 * 8.806744e-31 = -504442300000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011010100111111010111000010011;
		b = 32'b00011111110111001111111011101101;
		correct = 32'b11111010001110001111100011100000;
		#400 //-2.247296e+16 * 9.3595364e-20 = -2.401076e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010111000011010101100100000111;
		b = 32'b10111010111100100110110011001001;
		correct = 32'b10011011100101010100001101000111;
		#400 //4.5671925e-25 * -0.0018495555 = -2.469346e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010100010101011111000011101010;
		b = 32'b11111011011010110000100100001100;
		correct = 32'b10011000011010010000011000110000;
		#400 //3675479600000.0 * -1.22037325e+36 = -3.0117668e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010111110000100100011001110111;
		b = 32'b10111000100100010100100101100011;
		correct = 32'b10011110101010110010100011100111;
		#400 //1.2554744e-24 * -6.927808e-05 = -1.8122246e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111010000111010110111001101101;
		b = 32'b11001100000000100001011100011010;
		correct = 32'b10101101100110101110011011011101;
		#400 //0.00060055294 * -34102376.0 = -1.7610297e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101111111100011000011000100111;
		b = 32'b11000010001000000111000001111101;
		correct = 32'b11101101010000001011000010100111;
		#400 //1.49496135e+29 * -40.10985 = -3.7271676e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100100100010011011110111111000;
		b = 32'b00110010111010110110010110010010;
		correct = 32'b11110001000101011100110001001011;
		#400 //-2.032714e+22 * 2.740379e-08 = -7.417639e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100111010111010110111000111100;
		b = 32'b00001001011010000001010011011010;
		correct = 32'b11011101011101000100000001100000;
		#400 //-3.072967e-15 * 2.7935789e-33 = -1.1000108e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001101000101111001010111010011;
		b = 32'b01000100011101000110010100010000;
		correct = 32'b10001000000111101100100010001010;
		#400 //-4.671081e-31 * 977.5791 = -4.778213e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010110011011101001000111101011;
		b = 32'b11000001011001001101100100111010;
		correct = 32'b00010100100001010110111111111011;
		#400 //-1.927153e-25 * -14.303034 = 1.3473737e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110010000100101100010100101010;
		b = 32'b01100111101010110111011010100011;
		correct = 32'b01001001110110110010000111011010;
		#400 //2.9070828e+30 * 1.6194263e+24 = 1795131.2
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011011000110001111001011110000;
		b = 32'b00110110110000000001001110101001;
		correct = 32'b11100011110010111101100110110110;
		#400 //-4.305131e+16 * 5.7243346e-06 = -7.5207535e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110111000110001100001011111000;
		b = 32'b11010001110001110111100110111101;
		correct = 32'b11100100110001000000110010001000;
		#400 //3.0983733e+33 * -107092615000.0 = -2.8931718e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100000101100010011001011111001;
		b = 32'b10010001001000100111010101001100;
		correct = 32'b01001111000010111001110101000011;
		#400 //-3.0018697e-19 * -1.2815692e-28 = 2342339300.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010010000111001010011111100000;
		b = 32'b11110001100101111110010010100110;
		correct = 32'b10100000000001000000001101110000;
		#400 //168207840000.0 * -1.504277e+30 = -1.1181972e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110001001100001000100101100111;
		b = 32'b00011011011011001110001101010101;
		correct = 32'b01010101001111101100011110010100;
		#400 //2.5689475e-09 * 1.9594917e-22 = 13110274000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010000010011110001000100100000;
		b = 32'b00111100000000001110010011000111;
		correct = 32'b10010011110011011010000110011000;
		#400 //-4.0836744e-29 * 0.007867045 = -5.190862e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111100101100100100010101111001;
		b = 32'b01011001000001000000100010010101;
		correct = 32'b10100011001011001101001101001000;
		#400 //-0.021761643 * 2322758300000000.0 = -9.368879e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101010000111110101001101100000;
		b = 32'b00001000011100011000011010101011;
		correct = 32'b11100001001010001101111110100101;
		#400 //-1.4150963e-13 * 7.26816e-34 = -1.9469802e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101101010010010011110001110001;
		b = 32'b11101011000011101101110101110010;
		correct = 32'b01000001101101000100110000110000;
		#400 //-3.8924723e+27 * -1.7271321e+26 = 22.5372
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000110010010110000001110011100;
		b = 32'b10010010000001010110000101010101;
		correct = 32'b01110011110000101101001100110110;
		#400 //-12992.902 * -4.208737e-28 = 3.087126e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100111110001111110111111100011;
		b = 32'b00101101101110010010100100000100;
		correct = 32'b01111001100010100011011100010011;
		#400 //1.8883521e+24 * 2.105028e-11 = 8.970675e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110111001000011000100000011011;
		b = 32'b11001011110110101000100111100011;
		correct = 32'b11101010101111010011100010010110;
		#400 //3.2762513e+33 * -28644294.0 = -1.143771e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101110001101110101111000101100;
		b = 32'b00110000010111001000011101110101;
		correct = 32'b10111101010101001101110010001110;
		#400 //-4.1693024e-11 * 8.022803e-10 = -0.05196815
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011101101001000110001000000101;
		b = 32'b01000000000001010001001101010100;
		correct = 32'b00011101000111100001110100000011;
		#400 //4.351179e-21 * 2.0793047 = 2.0926125e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011000111010110010100010111100;
		b = 32'b11001001100010101100111010000010;
		correct = 32'b10001110110110001101100111011100;
		#400 //6.0787207e-24 * -1137104.2 = -5.3457902e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110111001000011010110001110000;
		b = 32'b00101000001000001111111001001111;
		correct = 32'b01001110100000001000101001110010;
		#400 //9.6364965e-06 * 8.936929e-15 = 1078278400.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101110111011100100101011101001;
		b = 32'b00111111000100000010101100111111;
		correct = 32'b11101111010100111001000101000101;
		#400 //-3.6873997e+28 * 0.5631599 = -6.5476957e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111111110100011100100110000111;
		b = 32'b11110011101011010000000110001110;
		correct = 32'b00001011100110110011011001111101;
		#400 //-1.6389626 * -2.7413907e+31 = 5.9785813e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101000101001001001101111101010;
		b = 32'b10111110000010001000000001011011;
		correct = 32'b11101010000110100101101101101010;
		#400 //6.2187537e+24 * -0.13330214 = -4.6651567e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011011001100010100010100111111;
		b = 32'b10000101010000011100110011010111;
		correct = 32'b01010101011010100010101001001000;
		#400 //-1.4663471e-22 * -9.1124395e-36 = 16091707000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101011110000011011100010101101;
		b = 32'b11000011110111000101110111110000;
		correct = 32'b00100111011000010000101111000000;
		#400 //-1.3764733e-12 * -440.7339 = 3.1231392e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000101000101101001101111110001;
		b = 32'b10010101000011001110010001010101;
		correct = 32'b01101111100010001101001111111101;
		#400 //-2409.7463 * -2.8452897e-26 = 8.469248e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110101001110111111001111110000;
		b = 32'b00110001001100001000001110010111;
		correct = 32'b01000011100010000100101110000001;
		#400 //7.0017904e-07 * 2.568617e-09 = 272.58987
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011101100110010100100110000110;
		b = 32'b10011000010111111010011011101010;
		correct = 32'b11000100101011110111010100111100;
		#400 //4.0574784e-21 * -2.8906345e-24 = -1403.6636
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000000000001101111101000101011;
		b = 32'b10001001100000111011101010101001;
		correct = 32'b01110110000000110010011111111000;
		#400 //-2.109019 * -3.1712637e-33 = 6.650406e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101101010111000101110111111100;
		b = 32'b00110100000111100010010101111011;
		correct = 32'b00111000101100100101110000101000;
		#400 //1.2526421e-11 * 1.4728532e-07 = 8.504867e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111001010101001000111010011110;
		b = 32'b11000001110110010111001000000000;
		correct = 32'b01110110111110100011111010111101;
		#400 //-6.897872e+34 * -27.180664 = 2.5377865e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010110101111111100110000110000;
		b = 32'b00111011011000010001010110001100;
		correct = 32'b00011010110110100010010000110110;
		#400 //3.0986575e-25 * 0.0034345118 = 9.022119e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011001000101101100100111010001;
		b = 32'b10000011110111001100101111001110;
		correct = 32'b01010100101011101101010010000100;
		#400 //-7.795575e-24 * -1.2977229e-36 = 6007118000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110001011100001110001010011000;
		b = 32'b01100010010100001001011001000100;
		correct = 32'b00001110100100111101000111100010;
		#400 //3.50534e-09 * 9.6193764e+20 = 3.6440408e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011000001001000011110001111100;
		b = 32'b10000101110101111010111101100100;
		correct = 32'b01010001110000101110111100111111;
		#400 //-2.122704e-24 * -2.0282931e-35 = 104654690000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110000100011111100010010000011;
		b = 32'b00111000011111000010011001101110;
		correct = 32'b00110111100100011111011001110100;
		#400 //1.0460471e-09 * 6.0117272e-05 = 1.740011e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011101100111010100000101100101;
		b = 32'b10110010011011010111010010110100;
		correct = 32'b01101010101010011000100101001100;
		#400 //-1.4164311e+18 * -1.3821751e-08 = 1.02478415e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010110001001110101110001100010;
		b = 32'b11001010000111111011010101111001;
		correct = 32'b10001011100001100010000111111100;
		#400 //1.3519303e-25 * -2616670.2 = -5.1666057e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010100010101111101111111100100;
		b = 32'b00100111111001010001111001011111;
		correct = 32'b10101011111100010011001110111011;
		#400 //-1.0898881e-26 * 6.3593197e-15 = -1.7138438e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111101100010011100110000100101;
		b = 32'b10101101101000100001100001111001;
		correct = 32'b11001111010110011010000000100101;
		#400 //0.067283906 * -1.8428136e-11 = -3651151000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001000100111111110011111010110;
		b = 32'b11001011010100001010100001110011;
		correct = 32'b00111100110001000010111110101111;
		#400 //-327486.7 * -13674611.0 = 0.023948519
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010110111100100011011000110000;
		b = 32'b11010000001101001001011100111000;
		correct = 32'b00000110001010111010110100010000;
		#400 //-3.9131406e-25 * -12119237000.0 = 3.2288672e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001101111111100010100110001100;
		b = 32'b11000101000100001110111101001000;
		correct = 32'b00001000011000000111011100001110;
		#400 //-1.5663961e-30 * -2318.955 = 6.7547496e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101111000101010000111100010111;
		b = 32'b11110011000001101001000000101011;
		correct = 32'b00111011100011011100100111101101;
		#400 //-4.613151e+28 * -1.0661192e+31 = 0.00432705
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010100100011100100010000001010;
		b = 32'b01010011000111001101110100100100;
		correct = 32'b00000000111010000010110100011000;
		#400 //1.4365172e-26 * 673725000000.0 = 2.1322012e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011011110100100000111110101010;
		b = 32'b10110100000010100110000100111000;
		correct = 32'b10100111010000100100110111111110;
		#400 //3.4751708e-22 * -1.288762e-07 = -2.6965188e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101110101000101000010100111110;
		b = 32'b11100011000010111010000011011011;
		correct = 32'b00001011000101001111110001010100;
		#400 //-7.3905757e-11 * -2.5756883e+21 = 2.8693594e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111100111001001010100110001;
		b = 32'b00110101000011101010001110100100;
		correct = 32'b11000010000011001000001100110100;
		#400 //-1.8666122e-05 * 5.313725e-07 = -35.128128
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111001011000011011100110110;
		b = 32'b11001011110011011011011000000010;
		correct = 32'b00101010110101100101000011111000;
		#400 //-1.0264854e-05 * -26962948.0 = 3.807022e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011110101101011010010011011101;
		b = 32'b01110000010111010100001000101000;
		correct = 32'b10101101110100100010101001010111;
		#400 //-6.5444147e+18 * 2.7390466e+29 = -2.3893039e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000101011111000111001011111111;
		b = 32'b01001100011000010010000101000101;
		correct = 32'b00111000100011111000100001011011;
		#400 //4039.1873 * 59016468.0 = 6.8441695e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111011100010111111000011000;
		b = 32'b01010110011001001100100110001010;
		correct = 32'b10100000100001110001101110110110;
		#400 //-1.4394078e-05 * 62888564000000.0 = -2.2888227e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111000110000100001000000000001;
		b = 32'b00011110110100111001000111101100;
		correct = 32'b01011001011010101101000011100000;
		#400 //9.253622e-05 * 2.2400846e-20 = 4130925300000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101100010101101110000101011110;
		b = 32'b01101100100010001001011111110101;
		correct = 32'b10111111010010010101110010001001;
		#400 //-1.0390976e+27 * 1.321052e+27 = -0.7865682
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000011010000010001011000001;
		b = 32'b00101101011110100100000100100110;
		correct = 32'b11000010011011010111011100011101;
		#400 //-8.4450497e-10 * 1.4225321e-11 = -59.36632
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001011110101011001001111010100;
		b = 32'b10110001000110111001010100010111;
		correct = 32'b10011010001011111011011010100011;
		#400 //8.226704e-32 * -2.2640216e-09 = -3.6336685e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001000010100001011001000110100;
		b = 32'b01101010001011001111101011011000;
		correct = 32'b00011101100110100110110111010001;
		#400 //213704.81 * 5.2279954e+25 = 4.087701e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101111110100000110010110010011;
		b = 32'b01001111101010100111011001111110;
		correct = 32'b00011111100111000111110000000101;
		#400 //3.7907152e-10 * 5719784400.0 = 6.627374e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011001100100011111010101110010;
		b = 32'b00101101101100011100111101100010;
		correct = 32'b10101011010100100010010001110111;
		#400 //-1.5091783e-23 * 2.0214667e-11 = -7.465759e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010001010000110011110001011010;
		b = 32'b10000010111011111001111110101101;
		correct = 32'b11001101110100001001010000010111;
		#400 //1.5401385e-28 * -3.5209543e-37 = -437420770.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110110100100001110110010000001;
		b = 32'b01010101001111100110010010001000;
		correct = 32'b00100000110000101101110011110001;
		#400 //4.319067e-06 * 13083687000000.0 = 3.3011085e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000110010110010000001100110100;
		b = 32'b01000110111101111010010011110110;
		correct = 32'b10111110111000000101010110101000;
		#400 //-13888.801 * 31698.48 = -0.4381535
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110110001101011010000000001000;
		b = 32'b00111101011010101011011010011111;
		correct = 32'b00111000010001100001100011011010;
		#400 //2.7064252e-06 * 0.057303067 = 4.7230023e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010000100010111011110000101100;
		b = 32'b00011001010101001010001001001101;
		correct = 32'b01110110101010000011101111001010;
		#400 //18754920000.0 * 1.09929195e-23 = 1.7060909e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110000010110100011100100000101;
		b = 32'b11010101000100010011110111101100;
		correct = 32'b10011010110000000101000100110011;
		#400 //7.938897e-10 * -9980946000000.0 = -7.9540523e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010101110000110011010110001111;
		b = 32'b00011110111110101010110110000001;
		correct = 32'b00110110010001110101101010010010;
		#400 //7.8844373e-26 * 2.6541539e-20 = 2.970603e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000011011001101001111110100110;
		b = 32'b00001001001001000011101111111000;
		correct = 32'b00111001101100111011111000000000;
		#400 //6.7774193e-37 * 1.976898e-33 = 0.00034283102
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010101010000111010101011010100;
		b = 32'b00101101010101101001100100101111;
		correct = 32'b11100111011010010110101010101000;
		#400 //-13446154000000.0 * 1.2198505e-11 = -1.10227885e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001111000110100110011001111110;
		b = 32'b01001010001011000100101111100011;
		correct = 32'b00000100011001010110100011101001;
		#400 //7.6125255e-30 * 2822904.8 = 2.6966993e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011000111100011111100010100110;
		b = 32'b01100101001011101011100111010101;
		correct = 32'b10110011001100010100001100101001;
		#400 //-2128401900000000.0 * 5.1569985e+22 = -4.1272106e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011111000101100011010111111100;
		b = 32'b00000111100001110011000110100100;
		correct = 32'b01010111000011100011011111001000;
		#400 //3.180839e-20 * 2.0341719e-34 = 156370230000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100111100101100010101001000110;
		b = 32'b01000001101101110111101110100010;
		correct = 32'b10100101010100011000001110100000;
		#400 //-4.1679196e-15 * 22.935368 = -1.8172457e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101111011010000001100001101011;
		b = 32'b10000100010010001100111001001011;
		correct = 32'b01101010100100111111000111101000;
		#400 //-2.1108952e-10 * -2.3604612e-36 = 8.942723e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100111001111000111011101011101;
		b = 32'b01001100000010100100011000001010;
		correct = 32'b11011010101011100111011010100010;
		#400 //-8.9000676e+23 * 36247590.0 = -2.4553542e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100110011010110110110101001001;
		b = 32'b01011010010111000110001101111100;
		correct = 32'b00001011100010001011101111101111;
		#400 //8.168011e-16 * 1.550847e+16 = 5.2668066e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001000001010011101111111110001;
		b = 32'b01011011010000010111101001110100;
		correct = 32'b10101100011000001100010011100001;
		#400 //-173951.77 * 5.445931e+16 = -3.1941604e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001011100110000110010011010010;
		b = 32'b00100100101011100000111000100000;
		correct = 32'b10100110011000000010001111111010;
		#400 //-5.869997e-32 * 7.54844e-17 = -7.776437e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000010010110011011101001010111;
		b = 32'b00010101111110101000010000100011;
		correct = 32'b01101011110111100111111001110110;
		#400 //54.431973 * 1.0118267e-25 = 5.3795745e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011101010011000101001011000110;
		b = 32'b01001110010011011011110101110000;
		correct = 32'b10001110011111100011110010111110;
		#400 //-2.7041968e-21 * 862936060.0 = -3.1337163e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010101111001011100110010100011;
		b = 32'b00111101100001100110111011100001;
		correct = 32'b10010111110110101100110101111000;
		#400 //-9.2815223e-26 * 0.06564117 = -1.4139787e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000101111000101010110010101100;
		b = 32'b10010111011111101100001100100111;
		correct = 32'b11101101111000111100011010010110;
		#400 //7253.584 * -8.2318143e-25 = -8.8116466e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011100100011001101001100101110;
		b = 32'b00010110111010011110111001111101;
		correct = 32'b11000101000110100001110000100100;
		#400 //-9.319012e-22 * 3.7793687e-25 = -2465.7588
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100101111001010001111001111101;
		b = 32'b01000011110011001000000011011100;
		correct = 32'b01100001100011110110100000111011;
		#400 //1.3524804e+23 * 409.0067 = 3.3067437e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100010011001001101011001001111;
		b = 32'b11111111000011111101000001111110;
		correct = 32'b00100010110010111010110001011100;
		#400 //-1.05532505e+21 * -1.9116216e+38 = 5.5205753e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011101001001011010101111110011;
		b = 32'b10010101010011101000010100001100;
		correct = 32'b01000111010011010101110101111010;
		#400 //-2.1926464e-21 * -4.1706324e-26 = 52573.477
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111100010110001010000110000110;
		b = 32'b00111101000001011100111001000100;
		correct = 32'b11111110110011110011101101000100;
		#400 //-4.4992488e+36 * 0.032667413 = -1.3772896e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011101111100110110010101011010;
		b = 32'b01010111111101001111100010101110;
		correct = 32'b10000101011111100101101010000100;
		#400 //-6.442636e-21 * 538697800000000.0 = -1.1959648e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001000011001101011110000111100;
		b = 32'b10111011100100101010110110000100;
		correct = 32'b00001100010010010101101010001100;
		#400 //-6.9434376e-34 * -0.004476251 = 1.5511725e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111001100100011010001010101001;
		b = 32'b01011101100011001101010010000100;
		correct = 32'b10011011100001000101111000010011;
		#400 //-0.00027777746 * 1.2684851e+18 = -2.1898362e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110100110010100101011110000;
		b = 32'b10110011010011011001101011101010;
		correct = 32'b11001010101111101101110110010101;
		#400 //0.29939985 * -4.7871175e-08 = -6254282.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101110010101110010010000100000;
		b = 32'b00101110100010100110000001010011;
		correct = 32'b00111111010001110000001000110001;
		#400 //4.8917426e-11 * 6.292624e-11 = 0.7773772
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100111111010011101011001111100;
		b = 32'b11011111010010111000110101011001;
		correct = 32'b10001000000100110000101101101011;
		#400 //6.4903036e-15 * -1.4667477e+19 = -4.4249625e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110010011101010101011000010100;
		b = 32'b01010000000110100100111010111100;
		correct = 32'b10100001110010111000001001101000;
		#400 //-1.4280449e-08 * 10355405000.0 = -1.3790333e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110000010001010100010011100101;
		b = 32'b00100000110000010011101011010110;
		correct = 32'b01001111000000101010110011111100;
		#400 //7.176609e-10 * 3.2734406e-19 = 2192374800.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001010100111000100001101011110;
		b = 32'b00101010011101110001101010111011;
		correct = 32'b11011111101000011110001101110110;
		#400 //-5120431.0 * 2.1947281e-13 = -2.3330594e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010011000000010111100100111111;
		b = 32'b00101000100110001011000000100010;
		correct = 32'b01101001110110010001010000000111;
		#400 //556084950000.0 * 1.6951775e-14 = 3.2803935e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001001101101110011011111100100;
		b = 32'b01000111010011110001010110010010;
		correct = 32'b10000001111000100111111100100100;
		#400 //-4.4108207e-33 * 53013.57 = -8.3201726e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000011011010011101101100101111;
		b = 32'b10001011011101001110110111101001;
		correct = 32'b01110111011101000110110100100101;
		#400 //-233.85619 * -4.7171674e-32 = 4.9575553e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010101100000101101101101010100;
		b = 32'b10111001010111100101101010101000;
		correct = 32'b00011011100101101010100001010101;
		#400 //-5.285262e-26 * -0.00021205342 = 2.49242e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110001100001011010010101101011;
		b = 32'b10110111110110100101011010111001;
		correct = 32'b00111001000111001011001011100011;
		#400 //-3.8896153e-09 * -2.6028009e-05 = 0.0001494396
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110100011011010010001110110111;
		b = 32'b11101010100110010011110000011001;
		correct = 32'b11001001010001100001011001011001;
		#400 //7.515251e+31 * -9.262473e+25 = -811365.56
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010000010010010101101111011010;
		b = 32'b00111110101010110101000100111101;
		correct = 32'b01010001000101100111001000001110;
		#400 //13512960000.0 * 0.33460417 = 40384913000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101011111110100101100100101011;
		b = 32'b00001111111110111110011001011010;
		correct = 32'b11011011011111100110110001011010;
		#400 //-1.7788317e-12 * 2.4839239e-29 = -7.161378e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000101011101011000111001011010;
		b = 32'b10010110010010110110010101101111;
		correct = 32'b10101110100110101000100000100001;
		#400 //1.15459905e-35 * -1.6430216e-25 = -7.0272906e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110011101011001001111100010011;
		b = 32'b10111000111101011110110010010010;
		correct = 32'b00111010001100111011000110100111;
		#400 //-8.0383096e-08 * -0.00011726575 = 0.00068547804
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001000100000100100111010010110;
		b = 32'b10100011100110100110000101100101;
		correct = 32'b11100100010110000001010010010100;
		#400 //266868.7 * -1.6737962e-17 = -1.5943918e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101100011010110010010010101110;
		b = 32'b10110100111111101111000110001101;
		correct = 32'b01110110111011000001111000100000;
		#400 //-1.1370831e+27 * -4.7486938e-07 = 2.3945177e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100101111110010111000111010101;
		b = 32'b00001001110000101111101010111000;
		correct = 32'b11011011101000111100000101011111;
		#400 //-4.327175e-16 * 4.6939576e-33 = -9.218607e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110101010011101100011001000101;
		b = 32'b11000111111010100011010100001110;
		correct = 32'b11101100111000100000001111000000;
		#400 //2.621178e+32 * -119914.11 = -2.1858796e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100101100110010010011001110110;
		b = 32'b10110010100000010110000001001000;
		correct = 32'b01110010100101111000010101110010;
		#400 //-9.040394e+22 * -1.506136e-08 = 6.002376e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011100100101100101011101001;
		b = 32'b11110011000100000110110101010110;
		correct = 32'b00011000000000100001100010110010;
		#400 //-19240402.0 * -1.1442693e+31 = 1.6814574e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011000100000100011110001011111;
		b = 32'b00101000110110100000001100011101;
		correct = 32'b01101111000110001110110111010000;
		#400 //1145566400000000.0 * 2.4204212e-14 = 4.732922e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011010010001110111110110001010;
		b = 32'b00011001110111010000000100111110;
		correct = 32'b00111111111001110001010000101101;
		#400 //4.1253645e-23 * 2.2851366e-23 = 1.8053032
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001101010101001010101011100000;
		b = 32'b01001100010000010000100001101011;
		correct = 32'b11000000100011010000010100001010;
		#400 //-222998020.0 * 50602412.0 = -4.406865
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111101011110110110010010111110;
		b = 32'b11001100111000011001101010010010;
		correct = 32'b11110000000011101010000111011010;
		#400 //2.0884957e+37 * -118281360.0 = -1.7657015e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001111011001001110101011000110;
		b = 32'b10001001000011110111100100111100;
		correct = 32'b11000101110011000011101001111100;
		#400 //1.12864836e-29 * -1.7270003e-33 = -6535.3105
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000111000010111100011011011011;
		b = 32'b01010101101010111000101011000010;
		correct = 32'b10110000110100001001100001100100;
		#400 //-35782.855 * 23576556000000.0 = -1.5177304e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011010001010101010011101101001;
		b = 32'b01110001101001101110110111100001;
		correct = 32'b10101000000000101101101100101001;
		#400 //-1.2008704e+16 * 1.6531869e+30 = -7.2639724e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000011001111000100011011110000;
		b = 32'b10110010001001111011011010111000;
		correct = 32'b01010000100011111011000110101110;
		#400 //-188.2771 * -9.762225e-09 = 19286290000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101011111010110000010010001111;
		b = 32'b00010110011100011001110001010001;
		correct = 32'b11010100111110010000001110111010;
		#400 //-1.669902e-12 * 1.951715e-25 = -8556075000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001110000011110101010011100101;
		b = 32'b10110010110111000010111001000101;
		correct = 32'b00011010101001101010011000100011;
		#400 //-1.7666986e-30 * -2.5632412e-08 = 6.89244e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001000001000001111100011011100;
		b = 32'b01000001101001011000001001000101;
		correct = 32'b11000101111110001111101110011000;
		#400 //-164835.44 * 20.688608 = -7967.449
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111011011000101111001100110000;
		b = 32'b01101000001001001010100111001000;
		correct = 32'b00010010101100000110101100010010;
		#400 //0.0034629814 * 3.1104e+24 = 1.1133556e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001110000010101011111101101100;
		b = 32'b00010100101101110100101001110011;
		correct = 32'b00111000110000011100100110001001;
		#400 //1.710198e-30 * 1.8507643e-26 = 9.240496e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111000110000011110001000000001;
		b = 32'b10101010111110101111110110010000;
		correct = 32'b01001101010001011100000010100110;
		#400 //-9.245054e-05 * -4.4584865e-13 = 207358560.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000111100010111011000110110100;
		b = 32'b00100111000101000010110010100001;
		correct = 32'b10011111111100010101100101001110;
		#400 //-2.101884e-34 * 2.056332e-15 = -1.0221521e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110000110011100101011100101110;
		b = 32'b00111011111001000100111100001111;
		correct = 32'b00110100011001110101111000000011;
		#400 //1.5013251e-09 * 0.0069674323 = 2.1547753e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101111100101000100100100010000;
		b = 32'b00110100100100010111000111010001;
		correct = 32'b11111010100000101000000000000101;
		#400 //-9.178422e+28 * 2.7091167e-07 = -3.3879757e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100110000100100101000100110100;
		b = 32'b01101011100100011110111110011100;
		correct = 32'b00111010000000000101010110011001;
		#400 //1.7274086e+23 * 3.5285153e+26 = 0.00048955675
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101110110101011001101101101101;
		b = 32'b00101000110010101000010111111000;
		correct = 32'b01000101100001110000000101011001;
		#400 //9.713728e-11 * 2.2484605e-14 = 4320.1685
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011000101110111100111110100011;
		b = 32'b01001001100010010010011000000001;
		correct = 32'b11001110101011110100100001111111;
		#400 //-1652003700000000.0 * 1123520.1 = -1470382000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110101000111010110000001000111;
		b = 32'b00111111011110111001111100111011;
		correct = 32'b01110101001000000001110101000010;
		#400 //1.9949789e+32 * 0.9828984 = 2.0296897e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001000000100101010111001100111;
		b = 32'b00100111001010101110010101111101;
		correct = 32'b11100000010110111011100111100000;
		#400 //-150201.61 * 2.3716645e-15 = -6.333173e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000001011011100110010101000110;
		b = 32'b00010000001101010001000011100000;
		correct = 32'b10110000101010001000011100011100;
		#400 //-4.3786356e-38 * 3.5708956e-29 = -1.2262009e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111111001010001100011011110100;
		b = 32'b01111001111010100011011110100001;
		correct = 32'b10000100101110000111100101001010;
		#400 //-0.6592858 * 1.5201572e+35 = -4.336958e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110100000110010001011110001101;
		b = 32'b11011110110010110111000111010010;
		correct = 32'b10010100110000001010001111010001;
		#400 //1.4257803e-07 * -7.3298646e+18 = -1.945166e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000101011111010011001000011110;
		b = 32'b01110100011001001011010110111011;
		correct = 32'b00010000100011011011010000101100;
		#400 //4051.1323 * 7.2481056e+31 = 5.589229e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001010000110011110010111101101;
		b = 32'b10101000110100001010001111110010;
		correct = 32'b10100000101111001101010011101011;
		#400 //7.409926e-33 * -2.3163739e-14 = -3.1989336e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111110100000011000100011101011;
		b = 32'b00111100010000011010010110001011;
		correct = 32'b11000001101010110011111010010101;
		#400 //-0.25299773 * 0.011819254 = -21.405558
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000100111010010100011010100111;
		b = 32'b10100110100011111011010011001110;
		correct = 32'b10011101110011111100011110111111;
		#400 //5.484292e-36 * -9.971625e-16 = -5.4998976e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001011011111000011110001011110;
		b = 32'b10001110011100100011100001010010;
		correct = 32'b10111100100001010100101011110101;
		#400 //4.857885e-32 * -2.985592e-30 = -0.016271094
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110100001111010111010010010110;
		b = 32'b01101111100010101010110001011100;
		correct = 32'b01000100001011101101111110100011;
		#400 //6.0040817e+31 * 8.58346e+28 = 699.4943
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000010001111101100110010111101;
		b = 32'b00011010110011000110001011011110;
		correct = 32'b11100110111011101111101110001001;
		#400 //-47.69994 * 8.453215e-23 = -5.642816e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000011100011101101011011111011;
		b = 32'b01011011000101000110010001011100;
		correct = 32'b00100111111101100110101111100101;
		#400 //285.67953 * 4.1768643e+16 = 6.8395695e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101111000001101011101001100001;
		b = 32'b10110101100010111011111000100111;
		correct = 32'b01111000111101101101000000110101;
		#400 //-4.169631e+28 * -1.0411649e-06 = 4.004775e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011010010001011000000101011100;
		b = 32'b00001101001100110100111100100001;
		correct = 32'b11001100100011001111110101001000;
		#400 //-4.084314e-23 * 5.525388e-31 = -73919040.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100011111011010010101101101111;
		b = 32'b11011110101100100001110111011101;
		correct = 32'b11000100101010100110111111110001;
		#400 //8.750016e+21 * -6.417329e+18 = -1363.4982
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100011011111100100001101110111;
		b = 32'b11000010000000000010111000011001;
		correct = 32'b10100000111111011110100000000110;
		#400 //1.3783654e-17 * -32.045017 = -4.3013407e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101111110111111100100000101001;
		b = 32'b11011100100011100001101100000100;
		correct = 32'b00010010110010011001000110101111;
		#400 //-4.0705686e-10 * -3.199932e+17 = 1.2720797e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101001000000110100010001011000;
		b = 32'b11111101110111101100110001001110;
		correct = 32'b10101010100101101101010000100110;
		#400 //9.918252e+24 * -3.7018678e+37 = -2.679256e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111001101111111000010100001000;
		b = 32'b11101111000001011100011001111011;
		correct = 32'b11001010001101110100000001011101;
		#400 //1.2430336e+35 * -4.1401454e+28 = -3002391.2
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001000100011100110001100001001;
		b = 32'b10101111110111001101110100111011;
		correct = 32'b10011000001001010000100111001010;
		#400 //8.569597e-34 * -4.017496e-10 = -2.1330692e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100110101011111110100000110;
		b = 32'b11001110101101000111101111000111;
		correct = 32'b10110101100101111100001100001001;
		#400 //1711.907 * -1514005400.0 = -1.1307139e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001100000010110101100101110001;
		b = 32'b10011111110100010011010010001110;
		correct = 32'b10101011101010101000010011010010;
		#400 //1.0735086e-31 * -8.860189e-20 = -1.2116092e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101110110101110000011010011111;
		b = 32'b11101111011110011000000101001100;
		correct = 32'b00111110110111001001111110001110;
		#400 //-3.327364e+28 * -7.721808e+28 = 0.4309048
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011010001110010100111101111101;
		b = 32'b00100110100101011110011010010101;
		correct = 32'b01110011000111100011110010000011;
		#400 //1.3040067e+16 * 1.0401451e-15 = 1.2536777e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010101101010000111100100100101;
		b = 32'b01000010111010011001001110000011;
		correct = 32'b01010010001110001010010110100001;
		#400 //23154783000000.0 * 116.78811 = 198263200000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010011111011100111101001110000;
		b = 32'b11000000011101100101100110101011;
		correct = 32'b00010010111101111101000111010101;
		#400 //-6.020038e-27 * -3.849223 = 1.5639619e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110000101110101110010100001101;
		b = 32'b01001010100011110100101101111001;
		correct = 32'b11100101101001101111001000111010;
		#400 //-4.6272894e+29 * 4695484.5 = -9.854764e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000111000000101101111000100010;
		b = 32'b11000010000101001110100000010000;
		correct = 32'b10000100011000001111110011011011;
		#400 //9.845392e-35 * -37.226624 = -2.6447179e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001111101100011011001101000010;
		b = 32'b10110110011001011010011101011100;
		correct = 32'b11011000110001100001011000010111;
		#400 //5962630000.0 * -3.4221075e-06 = -1742385400000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001100110110010000010000000111;
		b = 32'b10101100010000111001110000100010;
		correct = 32'b00100000000011100000000111011000;
		#400 //-3.3436568e-31 * -2.7797838e-12 = 1.2028478e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011000110000100010100100100000;
		b = 32'b00011101100010111111000001001001;
		correct = 32'b01111010101100011001100010011111;
		#400 //1707855100000000.0 * 3.7041443e-21 = 4.6106603e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110001110001010000111111011100;
		b = 32'b11100100100011101000001101110011;
		correct = 32'b00001100101100001111111001001001;
		#400 //-5.7352576e-09 * -2.1031277e+22 = 2.7270136e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000000000011001100010100100101;
		b = 32'b01001000111000110100010111000101;
		correct = 32'b00110110100111101001000001000110;
		#400 //2.1995327 * 465454.16 = 4.7255626e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010111010011110100000000001100;
		b = 32'b11001111010000100111101001110101;
		correct = 32'b11000111100010000110011111110011;
		#400 //227873990000000.0 * -3262805200.0 = -69839.9
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110100000010010000010110101111;
		b = 32'b11110111110001001100101000110010;
		correct = 32'b00111011101100100011111111011110;
		#400 //-4.342407e+31 * -7.982744e+33 = 0.0054397425
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000110100000001111101111001001;
		b = 32'b01100011010101111111110001100000;
		correct = 32'b10100010100110001110000100100000;
		#400 //-16509.893 * 3.9842355e+21 = -4.1438043e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010100001010111101000010001010;
		b = 32'b11001101001000011001000001110100;
		correct = 32'b11000110100010000001111011110010;
		#400 //2951752500000.0 * -169412420.0 = -17423.473
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110000101001101111111000011;
		b = 32'b11110011011100011000011011111001;
		correct = 32'b10001010000111011100101101111101;
		#400 //0.14538483 * -1.9135759e+31 = -7.597547e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011000100101101100100111110010;
		b = 32'b00101111000100110000110011110010;
		correct = 32'b10101001000000110100000100000101;
		#400 //-3.8978004e-24 * 1.3374171e-10 = -2.914424e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101010010000010010011000101001;
		b = 32'b10110011011110000110101010110000;
		correct = 32'b01110110010001110000101110010010;
		#400 //-5.8375722e+25 * -5.783903e-08 = 1.00927905e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100110101000000101101000100000;
		b = 32'b10110011011001111000100101011011;
		correct = 32'b01110010101100010100101101011100;
		#400 //-3.7862058e+23 * -5.3908803e-08 = 7.0233537e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101111110101000001110000010011;
		b = 32'b11011101100010100101001011100000;
		correct = 32'b01010001110001000100011101101010;
		#400 //-1.3128952e+29 * -1.2459094e+18 = 105376465000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110101101010000001001010011110;
		b = 32'b11100110001010000101101000111101;
		correct = 32'b10001110111111111001001100010111;
		#400 //1.2522394e-06 * -1.9875554e+23 = -6.3003996e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010010110100001010101000110010;
		b = 32'b11111100110011101100101101011000;
		correct = 32'b10010101100000010010100001100101;
		#400 //448104300000.0 * -8.5898996e+36 = -5.2166416e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010101110010011000111101010010;
		b = 32'b11001001110010111111110010110100;
		correct = 32'b11001011011111001111010000101101;
		#400 //27702174000000.0 * -1671062.5 = -16577581.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100101100100100111100000101011;
		b = 32'b01011011110011001111000110110011;
		correct = 32'b01001001001101101111010100111111;
		#400 //8.646028e+22 * 1.1537329e+17 = 749395.94
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100110000001001100101001001110;
		b = 32'b10010010111101010101100011011100;
		correct = 32'b11010010100010101000111001010100;
		#400 //4.6070874e-16 * -1.5483579e-27 = -297546680000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110010011011111011100010000110;
		b = 32'b10000000010010000111100011111111;
		correct = 32'b01110001110100111011001000001011;
		#400 //-1.3953587e-08 * -6.655561e-39 = 2.0965305e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101100001101011010110000011011;
		b = 32'b11010110011100000101001100010010;
		correct = 32'b10010101010000011000010110101010;
		#400 //2.5817185e-12 * -66059894000000.0 = -3.9081482e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100111111011000000000011001101;
		b = 32'b11001111001000000010011110011101;
		correct = 32'b11011000001111001001111010111110;
		#400 //2.2289865e+24 * -2686950700.0 = -829559900000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001010010111110110011111001010;
		b = 32'b00111010010111111010010101011110;
		correct = 32'b00001111011111111011100110000011;
		#400 //1.075658e-32 * 0.00085314165 = 1.2608199e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001111111111000011110111101101;
		b = 32'b01001101000010110001000001111111;
		correct = 32'b00000010011010000010110000110101;
		#400 //2.4872971e-29 * 145819630.0 = 1.7057355e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000100001010001001101011100011;
		b = 32'b01011000000000110111011010001011;
		correct = 32'b10101011101001000010100111011111;
		#400 //-674.4201 * 578180650000000.0 = -1.1664522e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110000101111111111110001010;
		b = 32'b00100101101011111110111010101001;
		correct = 32'b01010111110111010010110001100101;
		#400 //0.14843574 * 3.0519383e-16 = 486365500000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001000111100110000100111101100;
		b = 32'b11100101101010111100111100010000;
		correct = 32'b10100010101101010001000100111010;
		#400 //497743.38 * -1.0141804e+23 = -4.9078388e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011010000000011011010001000000;
		b = 32'b00101011011011000110111111010100;
		correct = 32'b10101110000011000110111110100000;
		#400 //-2.682218e-23 * 8.3999236e-13 = -3.1931457e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011100100000100110111100000100;
		b = 32'b00111110001010001011001101100101;
		correct = 32'b01011101110001011110111000110001;
		#400 //2.9371048e+17 * 0.16474684 = 1.7827989e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001000100010011001111110001100;
		b = 32'b00010001000001100110100010101001;
		correct = 32'b10110111000000110000111110100110;
		#400 //-8.282897e-34 * 1.0602987e-28 = -7.811852e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100010011100110000010101111001;
		b = 32'b10001100111110101101110111100101;
		correct = 32'b11010100111101111111111001111011;
		#400 //3.2935538e-18 * -3.8652147e-31 = -8521011000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000011001111001010101000101101;
		b = 32'b10101011101101111101100101010011;
		correct = 32'b01010111000000110101101001010111;
		#400 //-188.66475 * -1.3063252e-12 = 144424030000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010101001000000111100100100111;
		b = 32'b01111101000110011010001110000001;
		correct = 32'b00010111100001011011000110101100;
		#400 //11027638000000.0 * 1.2763803e+37 = 8.639774e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101101011100001001000000010011;
		b = 32'b10000110001010100010101101111100;
		correct = 32'b11100110101101001111001011100110;
		#400 //1.3674411e-11 * -3.2005394e-35 = -4.2725333e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110101001110100000111110001111;
		b = 32'b01000010100111100011011101001101;
		correct = 32'b00110010000101101000011011101000;
		#400 //6.931304e-07 * 79.10801 = 8.761823e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111110011000110011011100000101;
		b = 32'b10010101110111000010110111010000;
		correct = 32'b01101000000001000001011100100000;
		#400 //-0.22188957 * -8.892957e-26 = 2.4951158e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100101110001001101101000001000;
		b = 32'b01111011000000111111101110110100;
		correct = 32'b10101010001111101110100100100111;
		#400 //-1.16200725e+23 * 6.85296e+35 = -1.6956281e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011001011100001101001000110010;
		b = 32'b10101100010001001110110100110000;
		correct = 32'b01101100100111001000011111101101;
		#400 //-4236569200000000.0 * -2.798494e-12 = 1.5138746e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110100000011001000010111001110;
		b = 32'b11111011111010001101110011000001;
		correct = 32'b10110111100110100111110000111100;
		#400 //4.4533413e+31 * -2.4181806e+36 = -1.8416082e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011010100111110000010000101100;
		b = 32'b11001101100001101100000010000011;
		correct = 32'b11001100100101110000110001101010;
		#400 //2.2379554e+16 * -282595420.0 = -79192910.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011011110010111110111110110101;
		b = 32'b00001011110110111011000010101001;
		correct = 32'b11001111011011011010010001111101;
		#400 //-3.373844e-22 * 8.462154e-32 = -3986980000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101110110010011010001110101101;
		b = 32'b00000001011101001001000100011001;
		correct = 32'b01101100110100110001000011010110;
		#400 //9.1694964e-11 * 4.4919825e-38 = 2.0413028e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110000110011001011001011010010;
		b = 32'b00001001111000101110100101000100;
		correct = 32'b01100110011001101111000010010101;
		#400 //1.4893777e-09 * 5.4626883e-33 = 2.7264556e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100001010001001100001100110111;
		b = 32'b00101011101010110000110001110010;
		correct = 32'b01110101000100110011111000001110;
		#400 //2.2685178e+20 * 1.2153735e-12 = 1.8665192e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010001010101101111000111010001;
		b = 32'b10111100000000011011110100101011;
		correct = 32'b10010100110101000001000001001001;
		#400 //1.6956139e-28 * -0.007918636 = -2.1412953e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011100111100001010101100111010;
		b = 32'b11011010100101100010100111111010;
		correct = 32'b11000001110011010010010110000001;
		#400 //5.4193808e+17 * -2.11337e+16 = -25.643312
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011000110100011100100111101110;
		b = 32'b01110010100101111001010100100000;
		correct = 32'b00100101101100010010011010011011;
		#400 //1845321700000000.0 * 6.004802e+30 = 3.0730766e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111010001111111110100000111011;
		b = 32'b11001111110101111100010000100110;
		correct = 32'b10101001111000111011000100100100;
		#400 //0.0007320677 * -7239912400.0 = -1.0111554e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101010100001110101001101010010;
		b = 32'b11100000000101110101010001000001;
		correct = 32'b01001001111001001110110101010000;
		#400 //-8.179923e+25 * -4.361765e+19 = 1875370.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011011011101011001100001111001;
		b = 32'b00101111100110001101011101111111;
		correct = 32'b10101011010011011010110110100100;
		#400 //-2.0315192e-22 * 2.7801758e-10 = -7.3071605e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000000100101100101010001010001;
		b = 32'b00101010010010110101101101000101;
		correct = 32'b11010101101111010011111011011100;
		#400 //-4.6977925 * 1.8061687e-13 = -26009710000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011100001001101001001001110010;
		b = 32'b00110010001000110000100100000010;
		correct = 32'b00101001100000101100011011011101;
		#400 //5.511407e-22 * 9.489897e-09 = 5.807657e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000001111100011110010010101111;
		b = 32'b01000100101011100101001101110110;
		correct = 32'b00111100101100011001110010011001;
		#400 //30.236662 * 1394.6082 = 0.021681117
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011111111000111000111100010000;
		b = 32'b01010010111010110010010101001111;
		correct = 32'b10001100011101111011110110000001;
		#400 //-9.6374917e-20 * 504971620000.0 = -1.9085215e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001110100111101101100011100110;
		b = 32'b01000110110000111100101111001111;
		correct = 32'b00000111010011111011000010100100;
		#400 //3.9158873e-30 * 25061.904 = 1.5624859e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000101110000010011100111100111;
		b = 32'b00011111110010001001010010111010;
		correct = 32'b11100101011101101001110011110111;
		#400 //-6183.238 * 8.494934e-20 = -7.2787353e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100110101000101100111000011000;
		b = 32'b00111100010010100100100110000010;
		correct = 32'b00101001110011100000100011001001;
		#400 //1.129687e-15 * 0.012346627 = 9.149762e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100110111100101000011000110100;
		b = 32'b00101001111000001011000010101111;
		correct = 32'b11111100100010100010100011011011;
		#400 //-5.7264415e+23 * 9.978248e-14 = -5.738925e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000001000101011010111100001110;
		b = 32'b11100001001111110000010100101001;
		correct = 32'b00011111010010001001101000100111;
		#400 //-9.355238 * -2.2023125e+20 = 4.247916e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010001011001001001001111111000;
		b = 32'b00010001011011100110000001100010;
		correct = 32'b00111111011101010111101000100011;
		#400 //1.8031625e-28 * 1.880459e-28 = 0.9588949
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010011011000000101010100100001;
		b = 32'b00100101000111100110100011110001;
		correct = 32'b11101101101101010100010001111000;
		#400 //-963500900000.0 * 1.3739871e-16 = -7.012445e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110100001010100111000000100001;
		b = 32'b11000101100011110111100100101011;
		correct = 32'b00101110000110000000111001111110;
		#400 //-1.5873276e-07 * -4591.146 = 3.457367e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010101110101000111101110100101;
		b = 32'b01010101111111000101011101100100;
		correct = 32'b10111111010101111001000001010000;
		#400 //-29203440000000.0 * 34681534000000.0 = -0.8420458
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000011101100011011110000010100;
		b = 32'b01100011010011110111100111110110;
		correct = 32'b00011111110110110100110101101011;
		#400 //355.46936 * 3.8272642e+21 = 9.2878185e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010100001011100101010001111001;
		b = 32'b10010101011111101000100001111100;
		correct = 32'b01111110001011110101010110101010;
		#400 //-2994966000000.0 * -5.140256e-26 = 5.8264923e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100001111011001110010000100000;
		b = 32'b10001111000010100011000100010011;
		correct = 32'b01010010010110110110101110011000;
		#400 //-1.6052366e-18 * -6.813377e-30 = 235600740000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001101110001000101100100001100;
		b = 32'b11100111001101010010110100001110;
		correct = 32'b10100110000010101011100000000110;
		#400 //411771260.0 * -8.5557945e+23 = -4.8127766e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100001001001001000000001110010;
		b = 32'b00100101101101001100000100111011;
		correct = 32'b11111010111010001111101100100110;
		#400 //-1.896576e+20 * 3.135596e-16 = -6.048534e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111000110100101001110001011100;
		b = 32'b10011100110110000101110010110000;
		correct = 32'b01011011011110010011000111110000;
		#400 //-0.000100427045 * -1.431764e-21 = 7.0142176e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000100111101000001011111010001;
		b = 32'b00010010000100101011100001111010;
		correct = 32'b10110010010101001111001011000101;
		#400 //-5.7385996e-36 * 4.629686e-28 = -1.23952235e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101101110101110011011101000011;
		b = 32'b11011100001111111001100110110010;
		correct = 32'b00010001000011111100011011001001;
		#400 //-2.4467211e-11 * -2.1572284e+17 = 1.1341966e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100011010100101111011111110000;
		b = 32'b10011101010010010111110010101101;
		correct = 32'b01000101100001100000010111111100;
		#400 //-1.1436626e-17 * -2.6666584e-21 = 4288.748
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110010111101010110011010100101;
		b = 32'b00000001101000100001001101000111;
		correct = 32'b01110000110000011100111010010101;
		#400 //2.8568431e-08 * 5.9537063e-38 = 4.798428e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111101010000110101010001111101;
		b = 32'b11010110110101110111010100011010;
		correct = 32'b10100101111010000001010111010010;
		#400 //0.047687996 * -118448970000000.0 = -4.026037e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011111010100101101110101111011;
		b = 32'b11100011000000010000010110000000;
		correct = 32'b10111011110100010011001000011010;
		#400 //1.5194436e+19 * -2.3800263e+21 = -0.0063841464
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011111110001001011011100001001;
		b = 32'b00111100001100110011001000001011;
		correct = 32'b11100011000011001000001110100110;
		#400 //-2.8349616e+19 * 0.010937224 = -2.5920304e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110100000000011010001111101010;
		b = 32'b00000010101000011011000101001101;
		correct = 32'b11110000110011010100000011001111;
		#400 //-1.2073693e-07 * 2.375859e-37 = -5.081822e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111100111101000101111001011110;
		b = 32'b10011000110011011001010010010001;
		correct = 32'b11100011100110000010011010010010;
		#400 //0.029830154 * -5.314127e-24 = -5.613369e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111100100011101111111110001011;
		b = 32'b01010101110110110011010011110111;
		correct = 32'b10100110001001101111111111111110;
		#400 //-0.017455837 * 30127566000000.0 = -5.7939754e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011110010110011000011000001100;
		b = 32'b00111000100110001110011001001111;
		correct = 32'b00100101001101100001100110011001;
		#400 //1.15156046e-20 * 7.290823e-05 = 1.5794656e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011101000100111101011100101011;
		b = 32'b00001011110010000001111011010010;
		correct = 32'b01010000101111010001111100111011;
		#400 //1.9566527e-21 * 7.708357e-32 = 25383524000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001000100011100110100010010010;
		b = 32'b11100010011000011111010100011000;
		correct = 32'b00100101101000010101011110111001;
		#400 //-291652.56 * -1.0420446e+21 = 2.798849e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111001110001111111010001101011;
		b = 32'b11001101000001100111101101011010;
		correct = 32'b11101100001111100101000100110101;
		#400 //1.2977806e+35 * -141014430.0 = -9.203176e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010101000001101010111010110010;
		b = 32'b00101100010001011001111011000010;
		correct = 32'b11101000001011100111100000110011;
		#400 //-9255304000000.0 * 2.8083512e-12 = -3.2956362e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100010011110100011011110111101;
		b = 32'b10110101011000100110101000100010;
		correct = 32'b10101100100011010111010011101101;
		#400 //3.3910825e-18 * -8.4346004e-07 = -4.0204424e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110011101001001101101111100110;
		b = 32'b01011010001111011001011101000010;
		correct = 32'b00011000110111101001101011101011;
		#400 //7.6768444e-08 * 1.334127e+16 = 5.7542082e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110010101011101000010011100011;
		b = 32'b00001111101011110000100110010010;
		correct = 32'b01100010011111110011110111110010;
		#400 //2.0316696e-08 * 1.7260019e-29 = 1.17709584e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010010111011000100000001110101;
		b = 32'b10000111001000001001010001101011;
		correct = 32'b11001011001111000101000110101110;
		#400 //1.4909584e-27 * -1.2080678e-34 = -12341678.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110111011111010011011111110;
		b = 32'b01110001011100100001111010110010;
		correct = 32'b10000100111111010110010000010101;
		#400 //-7.1421955e-06 * 1.1989197e+30 = -5.9571925e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010100111010001010010100001111;
		b = 32'b10100010100111001100100001110000;
		correct = 32'b11110001101111011110111101001011;
		#400 //7993613000000.0 * -4.2496106e-18 = -1.8810225e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000110010010101110010111110110;
		b = 32'b10011000101101000011110111111111;
		correct = 32'b00101101000100000001011011100001;
		#400 //-3.8160926e-35 * -4.659151e-24 = 8.1905325e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001000100101001001001010101100;
		b = 32'b10010010110000000000100001011101;
		correct = 32'b11110101010001100001000001000101;
		#400 //304277.38 * -1.2118965e-27 = -2.5107538e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001101100100110011100100100000;
		b = 32'b10000011000101100111100110011111;
		correct = 32'b01001001111110100111011110110001;
		#400 //-9.073327e-31 * -4.4220652e-37 = 2051830.1
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110110011110011111100101010101;
		b = 32'b01101011010001111101011001100111;
		correct = 32'b11001010101000000001110100001001;
		#400 //-1.2675185e+33 * 2.4158872e+26 = -5246596.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000000011000001100001000100110;
		b = 32'b10010101001101100000010010111011;
		correct = 32'b10101010100010000001010111111110;
		#400 //8.885855e-39 * -3.675834e-26 = -2.4173713e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000100111110111111110100100010;
		b = 32'b00011000101001110010010011010101;
		correct = 32'b00101011110000001111100110010001;
		#400 //5.9242282e-36 * 4.320568e-24 = 1.3711689e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101101000101111110110011101110;
		b = 32'b00011011110110111001000101100101;
		correct = 32'b11010000101100010010001001001000;
		#400 //-8.635965e-12 * 3.632447e-22 = -23774511000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100001100011110000010011011011;
		b = 32'b00110110000100100000010001110101;
		correct = 32'b00101010111110101011111000111011;
		#400 //9.691342e-19 * 2.175829e-06 = 4.454092e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011000011111001101000011101001;
		b = 32'b00101000100110011111011110010000;
		correct = 32'b11101111010100100010110110000101;
		#400 //-1111896800000000.0 * 1.7093775e-14 = -6.504688e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110001100011000001001101000001;
		b = 32'b11111101100011001111110100001100;
		correct = 32'b10110011011111100101011101111101;
		#400 //1.3872377e+30 * -2.3425727e+37 = -5.9218554e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100001100000110011100000000101;
		b = 32'b11001101111110010011110100010110;
		correct = 32'b11010011000001101100011101001111;
		#400 //3.0257e+20 * -522691260.0 = -578869460000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100011110000010001110111001100;
		b = 32'b01000000000011110001100101100011;
		correct = 32'b10100011001011001011110101011001;
		#400 //-2.0937721e-17 * 2.2359245 = -9.364235e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010001000110000010111010110101;
		b = 32'b00010011001011101011100100111010;
		correct = 32'b11111101010111101111100100110011;
		#400 //-40851165000.0 * 2.2053211e-27 = -1.8523908e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101011000110101101011110011100;
		b = 32'b01001101111001111010001111011011;
		correct = 32'b00011100101010110010000000111010;
		#400 //5.501101e-13 * 485784420.0 = 1.1324161e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001010001010010010110010110011;
		b = 32'b11000100001111111010100000010011;
		correct = 32'b00000101011000011111100001101010;
		#400 //-8.145461e-33 * -766.62616 = 1.06250756e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001000010101110100110111001010;
		b = 32'b00111000010000010100011011011111;
		correct = 32'b00001111100011101001011001110010;
		#400 //6.479065e-34 * 4.608079e-05 = 1.406023e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001100001000000110010101010010;
		b = 32'b10001110111011110000111111100001;
		correct = 32'b01111100101010111100001010010111;
		#400 //-42046790.0 * -5.893334e-30 = 7.134636e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001111010101001000010011111000;
		b = 32'b11111101111010000011101111010011;
		correct = 32'b00010000111010100100010010101001;
		#400 //-3565484000.0 * -3.858644e+37 = 9.2402514e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001000000001101010001110111000;
		b = 32'b10100101101010001000001001101010;
		correct = 32'b11100001110011001000101101110101;
		#400 //137870.88 * -2.9231726e-16 = -4.716481e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010100110100010001110010100011;
		b = 32'b00110111010100100110001111011001;
		correct = 32'b00011100111111100111000111011011;
		#400 //2.1114902e-26 * 1.2540223e-05 = 1.6837741e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110000110110010001100111110100;
		b = 32'b01111000111001101111100001101111;
		correct = 32'b10110111011100001010000011000100;
		#400 //-5.3751698e+29 * 3.7477097e+34 = -1.4342546e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011010011010110100011010000001;
		b = 32'b01010101101110010110110000110000;
		correct = 32'b10000100001000100110101000000101;
		#400 //-4.8653814e-23 * 25484290000000.0 = -1.909169e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000101010000100011100100110000;
		b = 32'b10000110000111000111001001101001;
		correct = 32'b01111110100111101110100001010100;
		#400 //-3107.5742 * -2.9424394e-35 = 1.0561217e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100010111101010011000101000011;
		b = 32'b11110110111001010101011111101111;
		correct = 32'b10101011100010001101100001110100;
		#400 //2.261501e+21 * -2.3258193e+33 = -9.723459e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100110111011111101100101010000;
		b = 32'b11101000010111011011000010000101;
		correct = 32'b00111110000010100111110000100100;
		#400 //-5.6632715e+23 * -4.1875968e+24 = 0.13523918
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001111110100000110110101111010;
		b = 32'b11111100101001011011011000001011;
		correct = 32'b10010010101000001111111011011000;
		#400 //6993671000.0 * -6.88337e+36 = -1.0160243e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010011001100101010010111100;
		b = 32'b00010101011000011011011101100101;
		correct = 32'b11100100100000101001110111101011;
		#400 //-0.000878643 * 4.558306e-26 = -1.9275647e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110110110000100011110110101001;
		b = 32'b10000001110110111111000000000010;
		correct = 32'b11110100011000100001011100000101;
		#400 //5.7888287e-06 * -8.079229e-38 = -7.1650756e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111110010101101100101011100000;
		b = 32'b00011000010000101111011100010000;
		correct = 32'b11100101100011010000010001101001;
		#400 //-0.20975828 * 2.5198647e-24 = -8.324188e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110001111100011110001101111;
		b = 32'b01000101000010010101101000011001;
		correct = 32'b10110000101100010100100010001100;
		#400 //-2.8347383e-06 * 2197.631 = -1.2899064e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110101000110101000000100100;
		b = 32'b10111010010100100011111100110001;
		correct = 32'b11000011110001101101101001000111;
		#400 //0.3189708 * -0.00080202805 = -397.7053
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011010000100000000101101011011;
		b = 32'b00000110110101111101000000001110;
		correct = 32'b11010010101010101101111000001101;
		#400 //-2.9787675e-23 * 8.117972e-35 = -366934920000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000001100011110101110010111111;
		b = 32'b00000010010000011110001111011101;
		correct = 32'b01111110101111010100100101001110;
		#400 //17.920286 * 1.4244794e-37 = 1.2580236e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100101101001100010011100000100;
		b = 32'b11100010011111110101010100001101;
		correct = 32'b00000010101001101001011001000010;
		#400 //-2.8822848e-16 * -1.1775121e+21 = 2.4477752e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000110101111110110110111111111;
		b = 32'b01000010100010000101010001111100;
		correct = 32'b00000011101100111011101110100100;
		#400 //7.200784e-35 * 68.16501 = 1.0563755e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100000000010111110100001111100;
		b = 32'b10111001010111001000010010100110;
		correct = 32'b11100110001000100110101101101111;
		#400 //4.0325776e+19 * -0.0002103025 = -1.917513e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010011000011110110111001011111;
		b = 32'b01100010001011111100110011000010;
		correct = 32'b00110000010100001101110101011010;
		#400 //616032040000.0 * 8.1073364e+20 = 7.598452e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111100010011111100011110001001;
		b = 32'b11011101111110010100000000010011;
		correct = 32'b11011101110101010110011111110111;
		#400 //4.31541e+36 * -2.245047e+18 = -1.9221914e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101100000000101110111000011111;
		b = 32'b01100010011110011101001001011000;
		correct = 32'b00001001000001100010101100001111;
		#400 //1.8606295e-12 * 1.152099e+21 = 1.614991e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011000100110100101100110011100;
		b = 32'b10001010101000000001101110110111;
		correct = 32'b01001101011101101100101100000111;
		#400 //-3.989855e-24 * -1.5417865e-32 = 258781300.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110111011001111100011011010001;
		b = 32'b11110001101001000011000110111110;
		correct = 32'b01000101001101001010111101001100;
		#400 //-4.7009885e+33 * -1.6261016e+30 = 2890.956
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001111000111011010011011111101;
		b = 32'b11000011000101111011111100010101;
		correct = 32'b11001011100001001111101101010000;
		#400 //2644966700.0 * -151.74641 = -17430176.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101010000110010001111100001010;
		b = 32'b10010101100010011110010011010111;
		correct = 32'b01010100000011100010001010000001;
		#400 //-1.3599899e-13 * -5.5694905e-26 = 2441857000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001001001011011000001000111010;
		b = 32'b11010000110010100010001001010110;
		correct = 32'b00110111110110111011111100001110;
		#400 //-710691.6 * -27129983000.0 = 2.6195801e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001010100110010001101000001100;
		b = 32'b10011111000110010101000001110111;
		correct = 32'b01101010111111111010010100100010;
		#400 //-5016838.0 * -3.246557e-20 = 1.5452795e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110101110001101111111000101001;
		b = 32'b11001101101011001000010100101001;
		correct = 32'b10100111100100111010010000100101;
		#400 //1.482612e-06 * -361801000.0 = -4.097866e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100100110010100111001101110111;
		b = 32'b10000110000001110000011111110011;
		correct = 32'b01011110001111111110100011010001;
		#400 //-8.779914e-17 * -2.5396518e-35 = 3.457133e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111000101001010111111000110001;
		b = 32'b01100001001010110110111100001000;
		correct = 32'b10010110111101110010000011110011;
		#400 //-7.891318e-05 * 1.9764962e+20 = -3.9925796e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110010001010011100101110100010;
		b = 32'b11101000110110001111111100011001;
		correct = 32'b00001000110010000101000010011111;
		#400 //-9.883395e-09 * -8.197895e+24 = 1.2056016e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011101010010000100101100111111;
		b = 32'b11010010001010001101101101101011;
		correct = 32'b11001010100101111101010010001110;
		#400 //9.020437e+17 * -181308930000.0 = -4975175.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001110110110001110001110011100;
		b = 32'b00011000100001111000010111011110;
		correct = 32'b01110101110011001101100101111010;
		#400 //1819397600.0 * 3.5031853e-24 = 5.1935523e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100110111111101000110010110011;
		b = 32'b10010111000011100100101110111101;
		correct = 32'b01001111011001001111100111100010;
		#400 //-1.7662927e-15 * -4.597827e-25 = 3841581600.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010000010110000111111011101001;
		b = 32'b10101000000100111000000100100101;
		correct = 32'b01100111101110111101111001011011;
		#400 //-14528783000.0 * -8.188143e-15 = 1.7743685e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100011000000100100010111000011;
		b = 32'b11011100111110100110100101001011;
		correct = 32'b00000101100001010010111000010000;
		#400 //-7.062087e-18 * -5.6387612e+17 = 1.252418e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111101101011101011011011000101;
		b = 32'b01011110011101111010111101011001;
		correct = 32'b01011110101101001001010001001100;
		#400 //2.9029333e+37 * 4.4618954e+18 = 6.5060544e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110100010111100000000110011100;
		b = 32'b10011001001110000010001000101110;
		correct = 32'b11011010100110100101001111000010;
		#400 //2.0675947e-07 * -9.5194796e-24 = -2.171962e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001110011000001111101000011001;
		b = 32'b10001001010011111011011010101101;
		correct = 32'b01000100100010101010001101100101;
		#400 //-2.773055e-30 * -2.5002612e-33 = 1109.1061
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001110001111100100110010111010;
		b = 32'b00010110110001001011010011100000;
		correct = 32'b10110110111101111010100101110110;
		#400 //-2.345625e-30 * 3.1779656e-25 = -7.3809015e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101111001011111000000010100001;
		b = 32'b11010000001011100001011001000111;
		correct = 32'b10011110100000010000101001101101;
		#400 //1.5961855e-10 * -11682782000.0 = -1.3662718e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000011010001100110001111110011;
		b = 32'b00110001010001101010100010001000;
		correct = 32'b00010001011111111010011110011111;
		#400 //5.8301706e-37 * 2.890859e-09 = 2.0167605e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010010010111100101000011001111;
		b = 32'b00111111001001101111100000100001;
		correct = 32'b00010010101010100110110111010011;
		#400 //7.0150453e-28 * 0.65222365 = 1.0755582e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100010111010111011111101000011;
		b = 32'b01010110111101110000111001001001;
		correct = 32'b11001011011101000100100000101011;
		#400 //-2.1743834e+21 * 135820360000000.0 = -16009259.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011000000010001101000110010000;
		b = 32'b11110100100100101101010000000100;
		correct = 32'b10100010111011101000110001000110;
		#400 //601734600000000.0 * -9.306342e+31 = -6.465855e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010111101110001000111001101000;
		b = 32'b11101001110101111010010110100100;
		correct = 32'b00101101010110110001011101100101;
		#400 //-405843540000000.0 * -3.2587658e+25 = 1.2453903e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001100010001011111000101001110;
		b = 32'b11100000111001100000011011000010;
		correct = 32'b10101010110111000100101100011110;
		#400 //51889464.0 * -1.3260119e+20 = -3.9131973e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101100011001101010001001111110;
		b = 32'b01110010000110111010010101111111;
		correct = 32'b10111001101111011010101100101001;
		#400 //-1.11528114e+27 * 3.082896e+30 = -0.00036176413
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011001100100110111101000010001;
		b = 32'b01000001101111101011010111001100;
		correct = 32'b01010111010001011111011100111000;
		#400 //5188879400000000.0 * 23.838768 = 217665590000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101011010011110011000010000010;
		b = 32'b11011101000101101001011000001011;
		correct = 32'b00001101101100000001110100010010;
		#400 //-7.360849e-13 * -6.781795e+17 = 1.0853836e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111000100101011110110100001100;
		b = 32'b01110010000110111110101001101101;
		correct = 32'b11000101111101100010101001010011;
		#400 //-2.4326879e+34 * 3.088229e+30 = -7877.2905
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000010011011011110101111001001;
		b = 32'b10100101001000111101001011101100;
		correct = 32'b00011100101110011110010011100001;
		#400 //-1.7479677e-37 * -1.420946e-16 = 1.2301437e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000000100101001100111101100001;
		b = 32'b10000010100001100100001111001011;
		correct = 32'b00111101100011011101110111011000;
		#400 //-1.3666047e-38 * -1.9728442e-37 = 0.06927079
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011000001111011111101100001;
		b = 32'b00011001000011101101101100001000;
		correct = 32'b11110001011100110100001100100110;
		#400 //-8896353.0 * 7.385461e-24 = -1.20457656e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011010110101100110010101111001;
		b = 32'b11001011010101000001010001010111;
		correct = 32'b10001111000000010110010111111100;
		#400 //8.8672263e-23 * -13898839.0 = -6.3798325e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101001101000110000100110110111;
		b = 32'b01011011001000101000100000000101;
		correct = 32'b10001110000000000110011000100100;
		#400 //-7.2403394e-14 * 4.57485e+16 = -1.5826397e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010010100010111100100010101100;
		b = 32'b00110111111000000010000011010000;
		correct = 32'b11011010000111111010100101100001;
		#400 //-300183600000.0 * 2.671816e-05 = -1.1235189e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100001110001100111010000010001;
		b = 32'b10111110111101001100001111011010;
		correct = 32'b11100010010011111001000000000110;
		#400 //4.5760235e+20 * -0.47805673 = -9.572135e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000110111101011010110100001110;
		b = 32'b11010111000000110100011100001110;
		correct = 32'b10101111011011111000101011010100;
		#400 //31446.527 * -144341200000000.0 = -2.1786245e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001010101001001011101100000111;
		b = 32'b01101110011110111111010110000111;
		correct = 32'b00011011101001110101111101011101;
		#400 //5397891.5 * 1.949439e+28 = 2.768946e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010000101011000000101101011101;
		b = 32'b11111010111110001000010111101000;
		correct = 32'b00010101001100010011100001101101;
		#400 //-23091407000.0 * -6.452028e+35 = 3.5789377e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101000110001101011101011100101;
		b = 32'b11101001111000000110011001000100;
		correct = 32'b10111110011000101011011100111011;
		#400 //7.507809e+24 * -3.391029e+25 = -0.2214021
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100101010000010000001101001111;
		b = 32'b01110101011101101001011100101001;
		correct = 32'b00101111010010000110000011000110;
		#400 //5.696736e+22 * 3.1259056e+32 = 1.8224275e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100111010100111100100011101101;
		b = 32'b11000101000101101100111000011110;
		correct = 32'b11100001101100111100001000011010;
		#400 //1.00012575e+24 * -2412.8823 = -4.144942e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111101000000101011010010111110;
		b = 32'b00011100111111010010101111011001;
		correct = 32'b01011111100001000010101010011011;
		#400 //0.03191065 * 1.675347e-21 = 1.904719e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010001101101101011011110111100;
		b = 32'b11100000011100111001001000100101;
		correct = 32'b00110000110000000000101010100101;
		#400 //-98095825000.0 * -7.0204526e+19 = 1.3972864e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110100001001111001001111001110;
		b = 32'b11101011001100101011100110011110;
		correct = 32'b01001000011100000000100001001011;
		#400 //-5.3107386e+31 * -2.1606535e+26 = 245793.17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011010011000001000101100111101;
		b = 32'b11100000100001100001010111110110;
		correct = 32'b10111001010101100101101000111011;
		#400 //1.5800872e+16 * -7.729519e+19 = -0.00020442244
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110111001100001100001100000110;
		b = 32'b10110110111111110100110111100001;
		correct = 32'b10111111101100010011111001011001;
		#400 //1.0535825e-05 * -7.6086585e-06 = -1.3847152
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111101100110100010001110111;
		b = 32'b00011000001100001110110000111001;
		correct = 32'b01101111000000011011001001000011;
		#400 //91784.93 * 2.2866729e-24 = 4.013907e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111000011101100011000010010001;
		b = 32'b10001111100110111011001010111001;
		correct = 32'b01101000010010100110010010111001;
		#400 //-5.86962e-05 * -1.5353022e-29 = 3.823104e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000111100001110010101001010001;
		b = 32'b11000110010000101110100011111010;
		correct = 32'b01000000101100011000011110010111;
		#400 //-69204.63 * -12474.244 = 5.5478015
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011111110001101001011001111100;
		b = 32'b00101000100101010100110101000001;
		correct = 32'b10110110101010100100000100001110;
		#400 //-8.410522e-20 * 1.6575827e-14 = -5.073968e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000010000000000001101101011110;
		b = 32'b00101101010101001111110010110111;
		correct = 32'b11010100000110011111101001100111;
		#400 //-32.026726 * 1.2106919e-11 = -2645324200000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000101000011011011111111010111;
		b = 32'b00101111001100101100011010101001;
		correct = 32'b10010101010010101111101010110111;
		#400 //-6.6650236e-36 * 1.6259584e-10 = -4.0991354e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100101011001110110110000110;
		b = 32'b00011110001000110110010101100011;
		correct = 32'b01100110000001110111011110001001;
		#400 //1383.4226 * 8.6501144e-21 = 1.5993113e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101111101101000111000011100100;
		b = 32'b01010001000000100011001001111111;
		correct = 32'b11011110001100010110010101010011;
		#400 //-1.1168756e+29 * 34949560000.0 = -3.1956786e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000000001010100001111101100101;
		b = 32'b11000000110100101011010011101111;
		correct = 32'b10111110110011101011000100100100;
		#400 //2.6581662 * -6.5845866 = -0.40369523
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000100001110001000101101101001;
		b = 32'b11010000010010010001000110010111;
		correct = 32'b00110011011010101111011000100110;
		#400 //-738.1783 * -13493493000.0 = 5.470624e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110110101100100101110111010000;
		b = 32'b01010000110010000010011101011010;
		correct = 32'b11100101011001000010001000111100;
		#400 //-1.8088508e+33 * 26864177000.0 = -6.733319e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011000010111010000000101010101;
		b = 32'b00000011010100101101111000100001;
		correct = 32'b11010100100001100010011101010100;
		#400 //-2.8564253e-24 * 6.1968445e-37 = -4609483500000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010101101010000000001000011100;
		b = 32'b00010110000000101001011011010100;
		correct = 32'b01111111001001001010110101011011;
		#400 //23090877000000.0 * 1.0548909e-25 = 2.188935e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110100011011110110100000101110;
		b = 32'b10011001111111000011100001110111;
		correct = 32'b01011001111100101111111010010000;
		#400 //-2.229651e-07 * -2.6078995e-23 = 8549605000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101000111100110111111010101101;
		b = 32'b10001011111011111011111111010001;
		correct = 32'b01011100100000011111111111101101;
		#400 //-2.7033356e-14 * -9.2348065e-32 = 2.9273332e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011001110110010100110100110001;
		b = 32'b10110100101010100001110111000110;
		correct = 32'b01100100101000111000000011100000;
		#400 //-7645618000000000.0 * -3.168663e-07 = 2.4128846e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011001011110101100001100110111;
		b = 32'b10111000111101101001101001010100;
		correct = 32'b11100000000000100010100010111100;
		#400 //4411461600000000.0 * -0.0001175894 = -3.751581e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011100111111010000011010011100;
		b = 32'b01100100010010111111111001010101;
		correct = 32'b00111000000111101100010000110001;
		#400 //5.697635e+17 * 1.5052062e+22 = 3.7852853e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011101000100111101001111111011;
		b = 32'b01010101000011011001001110101010;
		correct = 32'b01000111100001011010011011011010;
		#400 //6.6575835e+17 * 9729084000000.0 = 68429.7
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101010101100111010011011001010;
		b = 32'b00110011000000000000101001000110;
		correct = 32'b10110111001100111001100001100000;
		#400 //-3.191252e-13 * 2.9811666e-08 = -1.0704709e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111011010010011010011110000001;
		b = 32'b00111101111100011111011100010101;
		correct = 32'b11111100110101010101100111011010;
		#400 //-1.04704905e+36 * 0.11814705 = -8.862253e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000000011000111011111010110111;
		b = 32'b00010100010110100010010010110000;
		correct = 32'b01101011100001011010001001001100;
		#400 //3.5585153 * 1.1013423e-26 = 3.2310712e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110000000110011111000011101100;
		b = 32'b00111101100110010001001111100001;
		correct = 32'b11110010000000001011100011010101;
		#400 //-1.9056985e+29 * 0.07474495 = -2.549602e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101100011101010111001110100011;
		b = 32'b11110101100000010010101100100001;
		correct = 32'b10110110011100110011101100111000;
		#400 //1.1869316e+27 * -3.27481e+32 = -3.6244292e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100000101011101100011010110001;
		b = 32'b11100100110001000110011111100011;
		correct = 32'b00111011011000111100111010110000;
		#400 //-1.0075158e+20 * -2.8984381e+22 = 0.0034760647
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010110101011011010000110001101;
		b = 32'b11000010011011010110000101110111;
		correct = 32'b11010011101110110100000000000011;
		#400 //95454680000000.0 * -59.34518 = -1608465600000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111010110010101011100011110100;
		b = 32'b00011111001110010100000100100110;
		correct = 32'b01011011000011000001000111000001;
		#400 //0.0015466497 * 3.9229163e-20 = 3.9426017e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100111000011100110011101100101;
		b = 32'b01011010011011001011010000100000;
		correct = 32'b01001100000110100000001101001001;
		#400 //6.724833e+23 * 1.6656536e+16 = 40373540.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001100011110010111000100101000;
		b = 32'b01101101010010101110011011100100;
		correct = 32'b00011110100111010101110000010011;
		#400 //65389730.0 * 3.9246939e+27 = 1.6661103e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011101000110100010110000110000;
		b = 32'b10001010010110100010010111010110;
		correct = 32'b01010010001101001110110010010000;
		#400 //-2.0404575e-21 * -1.0503434e-32 = 194265740000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100111001100000101011000010000;
		b = 32'b11001111101111101111111111010000;
		correct = 32'b00010110111011000101100011000111;
		#400 //-2.4471561e-15 * -6408872000.0 = 3.8183883e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000001111011010001001100011100;
		b = 32'b00100001000000010111000000000001;
		correct = 32'b01100000011010100111000100010101;
		#400 //29.63433 * 4.3855136e-19 = 6.7573227e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111010011101001110110110110101;
		b = 32'b01101101100111111111010000011001;
		correct = 32'b01001100010000111111111111110010;
		#400 //3.1793543e+35 * 6.1879016e+27 = 51380170.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101010000000010011100101011111;
		b = 32'b11100001110111011101110111000100;
		correct = 32'b01000111100101010001101011100001;
		#400 //-3.905559e+25 * -5.115888e+20 = 76341.76
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100110110111110110110011000111;
		b = 32'b10111110101110000111000011110111;
		correct = 32'b10100111100110110000110111011110;
		#400 //1.5503218e-15 * -0.36023685 = -4.3036177e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010010101010000000001111110101;
		b = 32'b00111111001110010111000010000100;
		correct = 32'b11010010111001111111001000101110;
		#400 //-360810450000.0 * 0.7243731 = -498100270000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010000100111100110100000111100;
		b = 32'b11011101011100011011010101001111;
		correct = 32'b10110010101001111100011000000011;
		#400 //21261050000.0 * -1.0885571e+18 = -1.9531404e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000010010010110100010000100110;
		b = 32'b00101101101001010001110110101011;
		correct = 32'b01010100000111011001001100011011;
		#400 //50.81655 * 1.8771503e-11 = 2707111500000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010111011011101111001000100011;
		b = 32'b01011100101000011111010111111101;
		correct = 32'b00111010001111001101011110100001;
		#400 //262723740000000.0 * 3.647035e+17 = 0.0007203762
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111011010001101100011000011100;
		b = 32'b01010011101001110011110000000101;
		correct = 32'b10100111000110000010001111011001;
		#400 //-0.0030330485 * 1436533000000.0 = -2.111367e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011011011100111101111011111101;
		b = 32'b00101101101110111010011110101011;
		correct = 32'b01101101001001100101100001011101;
		#400 //6.8643598e+16 * 2.1333898e-11 = 3.2175835e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111001100011010100011000000001;
		b = 32'b11101011010011101011011111001110;
		correct = 32'b10001101101011101111010000001111;
		#400 //0.00026945773 * -2.4990671e+26 = -1.0782333e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011111111011111011010001100101;
		b = 32'b11110010111011101101001010001101;
		correct = 32'b10101100100000000111100100001011;
		#400 //3.4545083e+19 * -9.4607325e+30 = -3.6514173e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011110110010111001001110011101;
		b = 32'b01000000001110100011100000000011;
		correct = 32'b10011110000010111110111001011111;
		#400 //-2.1554512e-20 * 2.9096687 = -7.407893e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001001000001011110000100101000;
		b = 32'b00001101110110110101000010001011;
		correct = 32'b11111010100111000100011000100000;
		#400 //-548370.5 * 1.3516307e-30 = -4.057103e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010100101101110011001100110000;
		b = 32'b01110000100010000101111110111010;
		correct = 32'b10100011101010111111001101100001;
		#400 //-6294702400000.0 * 3.376455e+29 = -1.8642932e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011111011100001001110000101100;
		b = 32'b00111101001111010011101110111010;
		correct = 32'b10100001101000101100000001111110;
		#400 //-5.095116e-20 * 0.046199538 = -1.1028499e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011101001111010101100101000101;
		b = 32'b11001010100010100000111111101101;
		correct = 32'b01010010001011111000110001110100;
		#400 //-8.527508e+17 * -4524022.5 = 188493920000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100011101001111001100110101011;
		b = 32'b00000101001111011101110011001011;
		correct = 32'b01011101111000011111101110011110;
		#400 //1.8171257e-17 * 8.9272906e-36 = 2.0354728e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101001001000010101000000111010;
		b = 32'b01001110000010100011100100100111;
		correct = 32'b10011010100101010110000111100001;
		#400 //-3.5818767e-14 * 579750340.0 = -6.178309e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011001010000010010010111111;
		b = 32'b01111011100000110110000011100001;
		correct = 32'b10001111001000111101000111010111;
		#400 //-11019455.0 * 1.3643117e+36 = -8.076934e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100010001000111110111011111000;
		b = 32'b10011011100111010100110000000011;
		correct = 32'b01000110000001010110011010000110;
		#400 //-2.2217128e-18 * -2.6022593e-22 = 8537.631
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111000001111000001101011011001;
		b = 32'b11111111111010010011011100100000;
		correct = 32'b11111111111010010011011100100000;
		#400 //-4.4847697e-05 * nan = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010111100110011110100111101011;
		b = 32'b00100100001010111100011111111010;
		correct = 32'b11110010111001010101111101101101;
		#400 //-338459900000000.0 * 3.72491e-17 = -9.086391e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010010110011010010110000001110;
		b = 32'b00001100001000000100000010100011;
		correct = 32'b01000110001000111110000100001010;
		#400 //1.2948179e-27 * 1.2345403e-31 = 10488.26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000010011111000110000010000011;
		b = 32'b00010110101010010011110100000000;
		correct = 32'b00101011001111101110000101011100;
		#400 //1.8541734e-37 * 2.734192e-25 = 6.781431e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111110111111001100110101111010;
		b = 32'b00011110000010100101111000000101;
		correct = 32'b11100000011010011101110001111001;
		#400 //-0.49375516 * 7.325102e-21 = -6.7405908e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110001010110000110011111011111;
		b = 32'b10110101100111001000100110001101;
		correct = 32'b10111011001100001111010001000111;
		#400 //3.149118e-09 * -1.1662938e-06 = -0.002700107
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110111101011000011010111101000;
		b = 32'b00011100100000010110111011001010;
		correct = 32'b01011010101010100100110111100101;
		#400 //2.05291e-05 * 8.565142e-22 = 2.3968196e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001101111010000001111101100010;
		b = 32'b00111100011101011001111011111101;
		correct = 32'b11010000111100011110111001100000;
		#400 //-486796350.0 * 0.014991519 = -32471450000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111001110001011110110000110010;
		b = 32'b01010010111101011011011010111101;
		correct = 32'b01100110010011100011010101001010;
		#400 //1.2845914e+35 * 527666400000.0 = 2.4344763e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100000101110101010101110000100;
		b = 32'b01101101111101101101101011000010;
		correct = 32'b10110010010000011001010111110011;
		#400 //-1.0760792e+20 * 9.549722e+27 = -1.1268173e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000110011010011001101100110000;
		b = 32'b01011110110011011001110011001110;
		correct = 32'b10100111000100010110110101001010;
		#400 //-14950.797 * 7.4079717e+18 = -2.0182038e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110010110100110101100111111100;
		b = 32'b11101111001101000101100000111111;
		correct = 32'b10000011000101100000000111010011;
		#400 //2.4604553e-08 * -5.5813985e+28 = -4.4083132e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000101010111110011100110100111;
		b = 32'b10110101011000110110010000010110;
		correct = 32'b10001111011110110100111101100101;
		#400 //1.0495999e-35 * -8.4709734e-07 = -1.2390546e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001111010110010010011110001100;
		b = 32'b11100100011110110101001011010111;
		correct = 32'b00101010010111010011000111110010;
		#400 //-3643247600.0 * -1.8544408e+22 = 1.9646071e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110010111011011100110110010000;
		b = 32'b11110111011101001100010101011110;
		correct = 32'b10111010111110001011011001011101;
		#400 //9.4203465e+30 * -4.964545e+33 = -0.0018975247
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111011011100111100101100000000;
		b = 32'b01111101001101010000111001111011;
		correct = 32'b00111101101011000101101000101011;
		#400 //1.2658455e+36 * 1.5041591e+37 = 0.08415636
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100000011111010101111010000010;
		b = 32'b11010000011011011101001011010100;
		correct = 32'b00001111100010000101110111101100;
		#400 //-2.1461204e-19 * -15960068000.0 = 1.3446813e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011110100110111001101011000001;
		b = 32'b00101011000101000110001011100101;
		correct = 32'b00110011000001100011100111111101;
		#400 //1.6475268e-20 * 5.2717406e-13 = 3.1252046e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010111101001110000110010110010;
		b = 32'b10111001110111010100000011001111;
		correct = 32'b10011101010000010100100010110100;
		#400 //1.0795327e-24 * -0.0004220069 = -2.5580924e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110110001101101110110101011011;
		b = 32'b00011000101110011111110001000101;
		correct = 32'b01011100111110111100101001011011;
		#400 //2.7258272e-06 * 4.8076106e-24 = 5.669817e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001100101001011110110110001001;
		b = 32'b00110011100101111111111010000001;
		correct = 32'b01011000100010111011101111101110;
		#400 //86993990.0 * 7.0777794e-08 = 1229114100000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010011000001100100001001111001;
		b = 32'b01110100000101111001100011010111;
		correct = 32'b10011110011000101011100011111100;
		#400 //-576640840000.0 * 4.8043017e+31 = -1.2002594e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110111001000100011101101110;
		b = 32'b00100111010111110111001010001010;
		correct = 32'b01010111000000101100010010001011;
		#400 //0.44585747 * 3.1009559e-15 = 143780660000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101001101001101100110100000011;
		b = 32'b00110111111001011101110111110101;
		correct = 32'b11110001001110011100001110010100;
		#400 //-2.5206228e+25 * 2.7402284e-05 = -9.1985866e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001000100110010010001000101101;
		b = 32'b10101100110111001010101111001110;
		correct = 32'b11011011001100011010011001011000;
		#400 //313617.4 * -6.2718502e-12 = -5.0003968e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101100111011111011000011110001;
		b = 32'b11100111111111000010101000101000;
		correct = 32'b11000100011100110101011000111000;
		#400 //2.3181508e+27 * -2.381628e+24 = -973.34717
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011101110100010110101110011111;
		b = 32'b10111100010011101100011000111110;
		correct = 32'b01100001000000011010001101010010;
		#400 //-1.8862912e+18 * -0.012620507 = 1.494624e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000000101110110100010001111101;
		b = 32'b10010011011101101101000000000010;
		correct = 32'b00101100110000100011110100001100;
		#400 //-1.7197807e-38 * -3.1152121e-27 = 5.520589e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100101010110100110100111001110;
		b = 32'b00011111110100111100001001011001;
		correct = 32'b01000101000001000000010110101100;
		#400 //1.8944334e-16 * 8.96835e-20 = 2112.3545
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100100011100100011000011110111;
		b = 32'b01000011110000000010100010100000;
		correct = 32'b00100000001000010101001111010111;
		#400 //5.251686e-17 * 384.31738 = 1.3664971e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010111111000010100101000101111;
		b = 32'b00010010010010000111111010101111;
		correct = 32'b01000101000011111101010001100000;
		#400 //1.4559011e-24 * 6.326502e-28 = 2301.2734
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000011110001000100111011011000;
		b = 32'b00100100101010011010100110011100;
		correct = 32'b01011110100101000001101000110100;
		#400 //392.61597 * 7.3579396e-17 = 5.3359497e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011011001111000101000101010001;
		b = 32'b11011110010101011011101100010000;
		correct = 32'b10111100011000011000111110011111;
		#400 //5.3006704e+16 * -3.8502302e+18 = -0.013767152
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001111101011101010000000000000;
		b = 32'b10111011101101111010010000110110;
		correct = 32'b01010011011100110110111001001110;
		#400 //-5859442700.0 * -0.0056042923 = 1045527660000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011111011100001101000011110011;
		b = 32'b11011100001011011110101110011110;
		correct = 32'b01000010101100010011101110110110;
		#400 //-1.7352637e+19 * -1.9581694e+17 = 88.61662
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000010101011110001111001001110;
		b = 32'b00011010010010011000111001001000;
		correct = 32'b10100111110111100110101111011100;
		#400 //-2.5731333e-37 * 4.168076e-23 = -6.173432e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000000001011110010011001101100;
		b = 32'b01010100010010101111111011001101;
		correct = 32'b00101011010111001110001001001111;
		#400 //2.73672 * 3487433000000.0 = 7.8473767e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111010100011001110011110000010;
		b = 32'b00001010100100000000110111010111;
		correct = 32'b01101111011110100110011100001111;
		#400 //0.0010750147 * 1.3871902e-32 = 7.7495843e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011111110011001001110111001100;
		b = 32'b10111000101000100011100100111001;
		correct = 32'b01100110101000010111001100001111;
		#400 //-2.948833e+19 * -7.7354205e-05 = 3.8121173e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001000001100111010110000001000;
		b = 32'b00011010001100000110100100000011;
		correct = 32'b10101101100000100101110111100000;
		#400 //-5.4068075e-34 * 3.6480775e-23 = -1.4820978e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010100000011101110111111010111;
		b = 32'b10010010101111111111010001101110;
		correct = 32'b11000000101111101010000010011011;
		#400 //7.216468e-27 * -1.2114051e-27 = -5.957105
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101010101111110111100100111001;
		b = 32'b10001001110101010010011100001101;
		correct = 32'b01100000011001011111011010001111;
		#400 //-3.401253e-13 * -5.1314608e-33 = 6.6282356e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010000000110101101100001011010;
		b = 32'b00010011000111110011001111000010;
		correct = 32'b10111100011110001111111001101000;
		#400 //-3.0537816e-29 * 2.009414e-27 = -0.015197374
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101011001110011110100011001110;
		b = 32'b01011010000010000001110010010000;
		correct = 32'b11010000101011101101010010000011;
		#400 //-2.2475067e+26 * 9578000000000000.0 = -23465302000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111111001101110010001000111100;
		b = 32'b11110000000010100001011010111100;
		correct = 32'b00001110101010011100000100000001;
		#400 //-0.7153661 * -1.7094566e+29 = 4.1847573e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100101111010101011011000111011;
		b = 32'b11010110110110000010110010110000;
		correct = 32'b11001110100010101111100111100111;
		#400 //1.3854941e+23 * -118843220000000.0 = -1165816700.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100000110101001000001000101101;
		b = 32'b01101000101111100110101100101001;
		correct = 32'b00110111100011101101100101010010;
		#400 //1.2250281e+20 * 7.193811e+24 = 1.7028917e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100111000000100101010111001101;
		b = 32'b01110000101001011000011000010000;
		correct = 32'b10110101110010011001001111000100;
		#400 //-6.154904e+23 * 4.098168e+29 = -1.5018672e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010001010011010001000000100011;
		b = 32'b00101100011010011000000111110000;
		correct = 32'b01100100011000001101000011001001;
		#400 //55046190000.0 * 3.3183421e-12 = 1.6588461e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111000011000101111000000011110;
		b = 32'b01110110010001000100001000010110;
		correct = 32'b11000001100101000000001001101011;
		#400 //-1.8411394e+34 * 9.95147e+32 = -18.50118
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010111000111001010001001001011;
		b = 32'b01110111111100010100010101111100;
		correct = 32'b00011110101001100011001000011111;
		#400 //172220860000000.0 * 9.7871317e+33 = 1.7596663e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100110010010000010011010100010;
		b = 32'b00000000111011100010000111101000;
		correct = 32'b11100100110101110010101100101011;
		#400 //-6.9441296e-16 * 2.1869011e-38 = -3.1753284e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010010101001010110110010101001;
		b = 32'b00010011010001001001011010010001;
		correct = 32'b00111110110101110110101100001101;
		#400 //1.0439751e-27 * 2.4812913e-27 = 0.4207386
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001111000001000010001010100111;
		b = 32'b00011110110000100000000100110110;
		correct = 32'b10101111101011100101110000100101;
		#400 //-6.514776e-30 * 2.054105e-20 = -3.1715888e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000001100000100110111010101010;
		b = 32'b10110101101101011010110011111000;
		correct = 32'b01001011001101111100101011110000;
		#400 //-16.304035 * -1.3535891e-06 = 12045040.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000101000111010001100010000011;
		b = 32'b01101110011010010011010001000100;
		correct = 32'b00010110001011000111001110110011;
		#400 //2513.532 * 1.8043298e+28 = 1.3930558e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101111111001110011000001110010;
		b = 32'b01110101110000000000101000111011;
		correct = 32'b00111001100110100001100000010110;
		#400 //1.4309921e+29 * 4.8687915e+32 = 0.00029391114
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110101010001100011110011101000;
		b = 32'b11101110100111011111111011011101;
		correct = 32'b11000110001000001001101000110010;
		#400 //2.5129641e+32 * -2.4448629e+28 = -10278.549
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100100100010011001011011010111;
		b = 32'b11011010010010010101111010000110;
		correct = 32'b10001001101011101110101010101100;
		#400 //5.966981e-17 * -1.41701e+16 = -4.210966e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111101011011011000010000011010;
		b = 32'b10001101001101101010110000110110;
		correct = 32'b11101111101001100110110111011001;
		#400 //0.05798731 * -5.629037e-31 = -1.0301462e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101000011111100101110000000100;
		b = 32'b00011100111010110110010001111100;
		correct = 32'b01001011000010100101000001001110;
		#400 //1.4119785e-14 * 1.557697e-21 = 9064526.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001001011111011011010101010010;
		b = 32'b10101101111111101100100011000010;
		correct = 32'b11011010111111101110101101000000;
		#400 //1039189.1 * -2.8965611e-11 = -3.5876652e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100101000110010011100000011101;
		b = 32'b11010100010110001110010011110001;
		correct = 32'b10010000001101001101100000101001;
		#400 //1.3289647e-16 * -3726215700000.0 = -3.5665264e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011110001100111001000001110110;
		b = 32'b11101011010111001010100001111001;
		correct = 32'b00110010010100000101001100001011;
		#400 //-3.234743e+18 * -2.6675927e+26 = 1.2126075e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011010110000110101110011111011;
		b = 32'b11001110000111011000111110000101;
		correct = 32'b10001100000111101011010111010101;
		#400 //8.080033e-23 * -660857150.0 = -1.2226595e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001001010110100110001110011101;
		b = 32'b00011000011011110100110011000110;
		correct = 32'b10110000011010011010000101000010;
		#400 //-2.6287633e-33 * 3.0928787e-24 = -8.499407e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101010011000100100110111110100;
		b = 32'b10000010110111100110010100111101;
		correct = 32'b01100111000000100011111111110110;
		#400 //-2.0099878e-13 * -3.2678076e-37 = 6.150875e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100110000111111011110101011001;
		b = 32'b01101100100011001011100001110010;
		correct = 32'b10111001000100010100110011000111;
		#400 //-1.8858728e+23 * 1.360965e+27 = -0.0001385688
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010000000010100110111010010110;
		b = 32'b10100111011011101111010011111000;
		correct = 32'b01101000000101000100111000101011;
		#400 //-9290013000.0 * -3.3161933e-15 = 2.8014087e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100011000101111001111001011101;
		b = 32'b11001101010101010010001101110111;
		correct = 32'b01010101001101100001101111001110;
		#400 //-2.7968696e+21 * -223491950.0 = 12514409000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010001101010110110110101100001;
		b = 32'b10100000110010000101100001011100;
		correct = 32'b10110000010110110000110010000011;
		#400 //2.7046453e-28 * -3.393979e-19 = -7.9689516e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000101010111111000110100110100;
		b = 32'b00101100100010101001110000000111;
		correct = 32'b00011000010011100111000011000000;
		#400 //1.05113445e-35 * 3.9395184e-12 = 2.66818e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101010100110110100110010010001;
		b = 32'b01101000010100111001111011001111;
		correct = 32'b00000001101110111101111000001111;
		#400 //2.758666e-13 * 3.9973953e+24 = 6.901159e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111001010000100111111000011100;
		b = 32'b11111101000001011111010111111010;
		correct = 32'b00111011101110011101011010011010;
		#400 //-6.311646e+34 * -1.1129032e+37 = 0.0056713345
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001000011110010100100100001101;
		b = 32'b10011111010101110110110001101111;
		correct = 32'b10101000100101000001111010110100;
		#400 //7.5016583e-34 * -4.5617715e-20 = -1.6444616e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100010101111001011101100111101;
		b = 32'b01101111011110110011100000101110;
		correct = 32'b00110010110000000101001010100110;
		#400 //1.7407399e+21 * 7.7748655e+28 = 2.2389326e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101011010011100110111010100000;
		b = 32'b10110000110000010010110011110110;
		correct = 32'b01111010000010001100100010101101;
		#400 //-2.4956113e+26 * -1.4055377e-09 = 1.7755564e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000101101101001010100110110011;
		b = 32'b10011100110111100100011110000001;
		correct = 32'b11101000010100000001000111111000;
		#400 //5781.2124 * -1.4709211e-21 = -3.9303348e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011001001111011010101101110000;
		b = 32'b01011111011010010111010110111111;
		correct = 32'b00111001010011111111101101011100;
		#400 //3336704300000000.0 * 1.6822562e+19 = 0.00019834697
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010110010011001101001101110000;
		b = 32'b01010100000010100000001010000000;
		correct = 32'b11000001101111011111100001010100;
		#400 //-56302122000000.0 * 2370989700000.0 = -23.746254
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110111100011010011001010100101;
		b = 32'b11000100100000100100011110100011;
		correct = 32'b10110010100010101011101000011001;
		#400 //1.6832093e-05 * -1042.2386 = -1.6149942e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100010100111110011111000000001;
		b = 32'b11000100010110011101110000101000;
		correct = 32'b11011101101110110001111011000101;
		#400 //1.4687501e+21 * -871.43994 = -1.6854289e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111111010110111011010011000001;
		b = 32'b11111000000100100111100000000000;
		correct = 32'b11000110110000000000000010101001;
		#400 //2.9203946e+38 * -1.1882957e+34 = -24576.33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111100101101011000000011111101;
		b = 32'b10000000011110110111001101110011;
		correct = 32'b11111011101111000011000100101011;
		#400 //0.022156233 * -1.1337181e-38 = -1.9542981e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100001010001110100011101111100;
		b = 32'b10100100110000100111111011010100;
		correct = 32'b00111100000000110010010111110110;
		#400 //-6.751843e-19 * -8.4348944e-17 = 0.008004656
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100101001000000011000010100011;
		b = 32'b00111110011011101101011100101000;
		correct = 32'b01100110001010111011001011101001;
		#400 //4.727974e+22 * 0.23324263 = 2.0270624e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110010110001011100010001010001;
		b = 32'b11001010110100000110101011001100;
		correct = 32'b10100111011100101110101100001100;
		#400 //2.3023093e-08 * -6829414.0 = -3.3711666e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110101101010100010001011110011;
		b = 32'b00111001001100110010010111001110;
		correct = 32'b00111011111100110001111110001000;
		#400 //1.2676159e-06 * 0.00017084854 = 0.0074195303
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000001011011000001100100101100;
		b = 32'b00011100000110101001001101001011;
		correct = 32'b10100100110000111000000111010011;
		#400 //-4.3364414e-38 * 5.1144697e-22 = -8.47877e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101100000001000101000000100010;
		b = 32'b01001001111000010000000100110000;
		correct = 32'b11100001100101101000101000101010;
		#400 //-6.398265e+26 * 1843238.0 = -3.4712092e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101111010001110111001010011011;
		b = 32'b00011111100000101010100000011001;
		correct = 32'b11001111010000110110010001101111;
		#400 //-1.813966e-10 * 5.5335236e-20 = -3278139100.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000011001011100001110010011;
		b = 32'b00100011110101001001001011101110;
		correct = 32'b11001100000010100101100111010010;
		#400 //-8.358764e-10 * 2.3047313e-17 = -36267850.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101000100100011000010101100001;
		b = 32'b01101100111000010011011001110101;
		correct = 32'b00111011001001010110101000001000;
		#400 //5.4976284e+24 * 2.1781238e+27 = 0.0025240202
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000001111000100010001111011110;
		b = 32'b00100100101111110011110111001010;
		correct = 32'b01011100100101110101101110101110;
		#400 //28.267513 * 8.293772e-17 = 3.408282e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011011110101001011001010110100;
		b = 32'b01001100110110000000000111110001;
		correct = 32'b01001110011111000001001111100111;
		#400 //1.1973836e+17 * 113250184.0 = 1057290700.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100001101111110110000010101100;
		b = 32'b01010001011101101010110100010000;
		correct = 32'b01001111110001101001110010000101;
		#400 //4.4128676e+20 * 66216590000.0 = 6664293000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100101000111011001000000101011;
		b = 32'b00100010011010010101111100001011;
		correct = 32'b01000010001011001101011101011001;
		#400 //1.3666425e-16 * 3.1627704e-18 = 43.2103
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011111110111100011101101001011;
		b = 32'b10110111000111100110000001101101;
		correct = 32'b00101000001100111001101110001001;
		#400 //-9.411875e-20 * -9.439985e-06 = 9.970222e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100001011110000001010010111011;
		b = 32'b00111010010100101011010010110101;
		correct = 32'b11100110100101101011010001100111;
		#400 //-2.860179e+20 * 0.00080377917 = -3.558414e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010100010111110011011110110111;
		b = 32'b01000110101001111000000010000110;
		correct = 32'b10001101001010101001001110000000;
		#400 //-1.1269611e-26 * 21440.262 = -5.256284e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111000001111111110100110111010;
		b = 32'b11010100011101001001101111000101;
		correct = 32'b11100011010010001101100110111000;
		#400 //1.5569832e+34 * -4202341600000.0 = -3.705037e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100010110001100011011100010101;
		b = 32'b11101101111011111101100000110100;
		correct = 32'b00110100010100111001000100001001;
		#400 //-1.8282122e+21 * -9.2785364e+27 = 1.970367e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110010000111001001001101111111;
		b = 32'b01101010110010000010110011000000;
		correct = 32'b00000110110010000011111000010010;
		#400 //9.113932e-09 * 1.20998245e+26 = 7.532284e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001010011000011011001000000011;
		b = 32'b00010000110101101010011100110010;
		correct = 32'b00111001000001101001010110101001;
		#400 //1.0866836e-32 * 8.466572e-29 = 0.00012834989
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100001111001011110101100110000;
		b = 32'b01000110110111001000110000101110;
		correct = 32'b00011010100001010111000001010010;
		#400 //1.5579897e-18 * 28230.09 = 5.5188974e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001111111100000011101100100000;
		b = 32'b00010101100010010101110100101100;
		correct = 32'b10111001110111111101101011001100;
		#400 //-2.3688601e-29 * 5.548086e-26 = -0.0004269689
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011010010101001110111010010011;
		b = 32'b10001011101101010100111111011111;
		correct = 32'b11001110000101100101001010010101;
		#400 //4.403329e-23 * -6.983884e-32 = -630498600.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011110110011101010111010110011;
		b = 32'b00111100001110001111110010001100;
		correct = 32'b10100010000011110000001100100111;
		#400 //-2.1883352e-20 * 0.011290681 = -1.9381783e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001110111000110000101110011011;
		b = 32'b01010101000111011011000101100000;
		correct = 32'b10111001001110000100101100110000;
		#400 //-1904594300.0 * 10836572000000.0 = -0.00017575617
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111101101010000100011000110011;
		b = 32'b10011110100011101011010100010100;
		correct = 32'b11011110100101101110111010010110;
		#400 //0.082165144 * -1.5109727e-20 = -5.4378975e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011011100000000100011011101010;
		b = 32'b10011110100100011111100111010000;
		correct = 32'b01111100011000001111011000011000;
		#400 //-7.221354e+16 * -1.5455792e-20 = 4.6722635e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001101111000101110011110010100;
		b = 32'b11000111011100111110001011100000;
		correct = 32'b00000101111011100010110011000110;
		#400 //-1.3984076e-30 * -62434.875 = 2.239786e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110010100010111000011111000101;
		b = 32'b10111000111001101010100011100101;
		correct = 32'b01111001000110101101101111110001;
		#400 //-5.5273666e+30 * -0.00010998714 = 5.0254666e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111111111111011000011011001101;
		b = 32'b10011001110100001001101000111100;
		correct = 32'b11111111111111011000011011001101;
		#400 //nan * -2.156899e-23 = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100001101110000000101100111010;
		b = 32'b11100010011001110010101101011100;
		correct = 32'b10111110110010111101000000000101;
		#400 //4.2437623e+20 * -1.06608056e+21 = -0.39807144
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100000000110110110101101001110;
		b = 32'b10100110000111110111001000101001;
		correct = 32'b01111001011110011000100011100110;
		#400 //-4.4796523e+19 * -5.531892e-16 = 8.097866e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001101101011010001101011010000;
		b = 32'b10110011001100001101111010111000;
		correct = 32'b11011001111110101000110011011010;
		#400 //363026940.0 * -4.1180755e-08 = -8815451500000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011001110000011001001001000011;
		b = 32'b00110001111010101101011101100011;
		correct = 32'b11100111010100110000001011111100;
		#400 //-6810686000000000.0 * 6.834783e-09 = -9.964744e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100101000000000101010101111110;
		b = 32'b00001111100001011101100110111011;
		correct = 32'b11010100111101010111001011111011;
		#400 //-1.1131196e-16 * 1.319868e-29 = -8433568300000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100100010101110010111011100101;
		b = 32'b10000001101110111101010100000101;
		correct = 32'b11100010000100101010001101111111;
		#400 //4.6660415e-17 * -6.899862e-38 = -6.7625144e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101100000110100010010000111101;
		b = 32'b00010001101010110010110001010000;
		correct = 32'b01011001111001101000011100111101;
		#400 //2.1904833e-12 * 2.7006353e-28 = 8110992600000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011111000111011100110011101010;
		b = 32'b11111011011010100000111010100010;
		correct = 32'b00100011001011001001100000011111;
		#400 //-1.137072e+19 * -1.21529425e+36 = 9.3563516e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010000011001101101110011001100;
		b = 32'b10100101000010100111001110110100;
		correct = 32'b01101010110101010110111100101110;
		#400 //-15492919000.0 * -1.2008794e-16 = 1.2901312e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000011100101000110111010011101;
		b = 32'b01000001111111000001111111111001;
		correct = 32'b10000001000101101011011010100101;
		#400 //-8.724054e-37 * 31.515612 = -2.768169e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100110011010001111111111100110;
		b = 32'b00101111010111001101110001001100;
		correct = 32'b11110110100001110000100100000100;
		#400 //-2.7507738e+23 * 2.0087149e-10 = -1.3694198e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011011001000100010111010010100;
		b = 32'b10001101110010110011101100010000;
		correct = 32'b11001100110011000100101011110111;
		#400 //1.3415376e-22 * -1.252506e-30 = -107108280.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110110101111100110110110001000;
		b = 32'b01110111111111110111000000011111;
		correct = 32'b10111110001111101101100011001011;
		#400 //-1.9311679e+33 * 1.0361795e+34 = -0.18637387
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111110100100110011110111011100;
		b = 32'b11111001010001001011010101101100;
		correct = 32'b01000100101111111001111101101101;
		#400 //-9.785885e+37 * -6.3835616e+34 = 1532.982
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000001101000011110010111001011;
		b = 32'b11001110110000010000010000001111;
		correct = 32'b10110010010101101011101000110111;
		#400 //20.237204 * -1619134300.0 = -1.249878e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100111100110111101011010000100;
		b = 32'b10000011110010100001011111111101;
		correct = 32'b11100011010001010110011111110010;
		#400 //4.325372e-15 * -1.1878e-36 = -3.6414986e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000011111111000000100100110101;
		b = 32'b00000101010011001011100010100111;
		correct = 32'b01111110000111011001010101000010;
		#400 //504.07193 * 9.625949e-36 = 5.2365947e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101001010100011100011000111011;
		b = 32'b00000101101111101001100001101100;
		correct = 32'b11100011000011001110000101010100;
		#400 //-4.657926e-14 * 1.7923505e-35 = -2.5987808e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011111001010001100001011010000;
		b = 32'b10111010011011001100011000100011;
		correct = 32'b01100100001101100111011011100001;
		#400 //-1.2160511e+19 * -0.000903221 = 1.3463494e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101101100000011101010010011000;
		b = 32'b01011111011111101010010000111010;
		correct = 32'b11001101100000101000010111101000;
		#400 //-5.022572e+27 * 1.8348855e+19 = -273726720.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100011010111101100111010011100;
		b = 32'b01010010011001011000010001111100;
		correct = 32'b01010000011110001000001111101001;
		#400 //4.110065e+21 * 246442560000.0 = 16677578000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100001100010000011011101001111;
		b = 32'b01001101010111010011000010101100;
		correct = 32'b10010011100111011010011100110001;
		#400 //-9.230359e-19 * 231934660.0 = -3.9797235e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001011110001110001111100100000;
		b = 32'b00011111101100101001101100011001;
		correct = 32'b01101011100011101011001111101101;
		#400 //26099264.0 * 7.564252e-20 = 3.450343e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111001011000110101010100111;
		b = 32'b00010011100111101010100011111111;
		correct = 32'b01110011000010110001100100011110;
		#400 //44138.652 * 4.005145e-27 = 1.1020488e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011110111011111011010001011010;
		b = 32'b10111100101011101100001001101111;
		correct = 32'b10100001101011111001000101101000;
		#400 //2.5379701e-20 * -0.021332948 = -1.189695e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010111000011111101110101111110;
		b = 32'b00111011001111100101101100010010;
		correct = 32'b11011011010000010111101000101000;
		#400 //-158181460000000.0 * 0.0029045981 = -5.4458983e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111001101010010111110011111;
		b = 32'b00011011110110101001100100010011;
		correct = 32'b01101010110101000010111111011001;
		#400 //46383.62 * 3.6163997e-22 = 1.2825911e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001101101011100101001101100101;
		b = 32'b11001011001101101000000100110011;
		correct = 32'b01000001111101001000011100000011;
		#400 //-365587620.0 * -11960627.0 = 30.565924
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110100100110110000100110101000;
		b = 32'b00100010000111010000010010001011;
		correct = 32'b11010001111111001100010110010100;
		#400 //-2.8878026e-07 * 2.1279873e-18 = -135705820000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110000000100101011000011110001;
		b = 32'b01101110000110011001000011111100;
		correct = 32'b00000001011101001000100111110100;
		#400 //5.336594e-10 * 1.188162e+28 = 4.49147e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100011001011100111110110011010;
		b = 32'b01100111010110110001100101000111;
		correct = 32'b00111011010010111110000011111101;
		#400 //3.218784e+21 * 1.03466454e+24 = 0.0031109445
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001111101010100101100100001010;
		b = 32'b01011101101111101111101011111100;
		correct = 32'b10110001011001000101011111001111;
		#400 //-5715924000.0 * 1.7201986e+18 = -3.322828e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111000110111111111011110001111;
		b = 32'b11010011010001101011100011011000;
		correct = 32'b00100101000100000100001010111101;
		#400 //-0.0001067958 * -853504700000.0 = 1.2512621e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000111010100101011001011100011;
		b = 32'b10000010011100011110111010110111;
		correct = 32'b01000100010111101111001100111110;
		#400 //-1.5851214e-34 * -1.7774391e-37 = 891.80066
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010111110101111001001100010111;
		b = 32'b10100110110101011010000100100001;
		correct = 32'b11110000100000010010101001011101;
		#400 //474053500000000.0 * -1.4823518e-15 = -3.1979824e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010101001100001010111011000110;
		b = 32'b10110101111001001000000010011101;
		correct = 32'b00011110110001011111000111000101;
		#400 //-3.568079e-26 * -1.7024755e-06 = 2.095818e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010111010101010100011000000110;
		b = 32'b11001011011000000100110111101001;
		correct = 32'b01001011011100110110100100010100;
		#400 //-234496730000000.0 * -14700009.0 = 15952148.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100100001011011111010101111101;
		b = 32'b01000001010101110000111111100100;
		correct = 32'b11100010010011110001001010011110;
		#400 //-1.2835904e+22 * 13.44138 = -9.549544e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001111111101100110011110001011;
		b = 32'b10010111110101011110100010111000;
		correct = 32'b01110111100100110111000111011100;
		#400 //-8267962000.0 * -1.3823549e-24 = 5.98107e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110101010001001000001110011011;
		b = 32'b01001100111011000011111101010110;
		correct = 32'b01100111110101001111000111010000;
		#400 //2.491112e+32 * 123861680.0 = 2.0112047e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111011011111110011001000111;
		b = 32'b10111010100011000011000100101101;
		correct = 32'b00111100010110110000100101000010;
		#400 //-1.4299126e-05 * -0.0010695808 = 0.013368906
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100001100000101010000001101111;
		b = 32'b11001011111111000010000001000100;
		correct = 32'b10010101000001001010001001000000;
		#400 //8.851609e-19 * -33046664.0 = -2.678518e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010100011010011010001000111000;
		b = 32'b00100001101000001010111111110000;
		correct = 32'b01110010001110100001101110001000;
		#400 //4013795800000.0 * 1.0888592e-18 = 3.6862397e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000111010110100101100000100101;
		b = 32'b01111101110110110101001011010000;
		correct = 32'b10001000111111101101101101101010;
		#400 //-55896.145 * 3.6441365e+37 = -1.5338653e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100111101100110010110000111111;
		b = 32'b11100000111101111100010111100100;
		correct = 32'b00000110001110010001111100111110;
		#400 //-4.973045e-15 * -1.4283142e+20 = 3.4817586e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110011101110110101110101001010;
		b = 32'b00000000100110101011001011011000;
		correct = 32'b01110010100110110000011100110111;
		#400 //8.724835e-08 * 1.4206823e-38 = 6.141299e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110011011011001110110000100100;
		b = 32'b01010000101100011110111101000101;
		correct = 32'b10100010001010100110111100001011;
		#400 //-5.51628e-08 * 23881984000.0 = -2.3098082e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001101000001111111111010101101;
		b = 32'b10101100010011010011000101001000;
		correct = 32'b10100000001010011010101100011010;
		#400 //4.190664e-31 * -2.9159609e-12 = -1.437147e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000101101101010100110101100100;
		b = 32'b11110000001111001011001101011001;
		correct = 32'b10010100111101011111011010010010;
		#400 //5801.674 * -2.336e+29 = -2.4835933e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011011001010111110111001000101;
		b = 32'b00100010000011011001011100111111;
		correct = 32'b11111000100110110110110101111110;
		#400 //-4.83942e+16 * 1.9189132e-18 = -2.5219587e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101011111101001100100011000011;
		b = 32'b01001001001000101001011101101111;
		correct = 32'b00100010010000001011010011000011;
		#400 //1.7392965e-12 * 665974.94 = 2.6116547e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011111100101001111101101011011;
		b = 32'b11011010110000000100100001010110;
		correct = 32'b00000100010001100101100110111111;
		#400 //-6.309627e-20 * -2.7061365e+16 = 2.3315998e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101110101001001100011100000000;
		b = 32'b10100011110100011000111010101001;
		correct = 32'b11001010010010010100101110111010;
		#400 //7.493206e-11 * -2.2720244e-17 = -3298030.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111101011101100000100011100;
		b = 32'b10000100111100010011100111111010;
		correct = 32'b01110010001110010111010011110110;
		#400 //-2.083234e-05 * -5.671207e-36 = 3.673352e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000000111011000010100110001101;
		b = 32'b11110101100101111011111111111110;
		correct = 32'b10001010110001110011001110000010;
		#400 //7.380072 * -3.8473188e+32 = -1.9182378e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010100011101101000100010110011;
		b = 32'b10111010111010111110101111000101;
		correct = 32'b11011001000001011100001000010101;
		#400 //4235421500000.0 * -0.0017999342 = -2353098000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000011111110001101011110001011;
		b = 32'b00011010100000101111101011110001;
		correct = 32'b01101000111100110010111000010011;
		#400 //497.68393 * 5.417216e-23 = 9.18708e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000111111100100001101010011111;
		b = 32'b01000110001001100001100001010000;
		correct = 32'b00000001001110101001001101101011;
		#400 //3.642776e-34 * 10630.078 = 3.4268572e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001000100010011010011000101100;
		b = 32'b00001111000001010101110101000000;
		correct = 32'b00111001000001000001110011001101;
		#400 //8.284454e-34 * 6.5753656e-30 = 0.0001259923
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110001111000000100101000001010;
		b = 32'b01011101100000100101100101000000;
		correct = 32'b11010011110111000011111101111010;
		#400 //-2.2212528e+30 * 1.1740761e+18 = -1891915500000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000010101000110110110001110111;
		b = 32'b10010100110000000110100011011000;
		correct = 32'b10101101010110010110111100111000;
		#400 //2.4012953e-37 * -1.9428399e-26 = -1.2359717e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101010100110101011100101011111;
		b = 32'b00100100110100111010001111100100;
		correct = 32'b01000101001110110010011110000000;
		#400 //2.7484522e-13 * 9.1784305e-17 = 2994.4688
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000101010011110000101010100001;
		b = 32'b00110001000100000001000111110100;
		correct = 32'b11010011101101111111001010000100;
		#400 //-3312.6643 * 2.0964963e-09 = -1580095500000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110101000001000100000110111101;
		b = 32'b11011101110101000001111001100100;
		correct = 32'b11010110100111111001110111101111;
		#400 //1.676554e+32 * -1.9105955e+18 = -87750334000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101000110010111011000101110110;
		b = 32'b00001100100000010000101000110100;
		correct = 32'b11011011110010100000110101000000;
		#400 //-2.2614489e-14 * 1.9881738e-31 = -1.1374503e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100101000011100100100011111100;
		b = 32'b00111100010011011001101100011011;
		correct = 32'b10101000001100010010100011000101;
		#400 //-1.2341265e-16 * 0.012549187 = -9.834314e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011101010001010110100111000101;
		b = 32'b11000000000100000011000101001110;
		correct = 32'b00011100101011110011111001110110;
		#400 //-2.6127414e-21 * -2.2530093 = 1.1596674e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101000010011110000001010101001;
		b = 32'b10110100101101100101111010001110;
		correct = 32'b01110011000100010100101101111100;
		#400 //-3.9103157e+24 * -3.396894e-07 = 1.1511445e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000100101101011010001111111011;
		b = 32'b00100100111000111110100010010001;
		correct = 32'b10011111010011000000011101111001;
		#400 //-4.2703488e-36 * 9.883954e-17 = -4.320486e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111000110100001011010100100001;
		b = 32'b11001011110100011000100001101010;
		correct = 32'b10101100011111101111110111011100;
		#400 //9.951951e-05 * -27463892.0 = -3.6236491e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100001000100110000101000000011;
		b = 32'b01011011000010100010110011011000;
		correct = 32'b00000101100010000011011000010001;
		#400 //4.981879e-19 * 3.8892853e+16 = 1.280924e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111110000111000100100010010;
		b = 32'b00010101100101000111100100110001;
		correct = 32'b11100001101010001001001010010000;
		#400 //-2.330964e-05 * 5.996793e-26 = -3.8870174e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001111000011010001111111100011;
		b = 32'b11000111000111010000011101101011;
		correct = 32'b00000111011001100001001001001100;
		#400 //-6.957978e-30 * -40199.418 = 1.7308654e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110010000110111111010100100100;
		b = 32'b11011011011010011100010001001100;
		correct = 32'b10010110001010101100101001011101;
		#400 //9.077926e-09 * -6.57995e+16 = -1.3796345e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111101101100110101100011010000;
		b = 32'b01100001111100011101011111111101;
		correct = 32'b01011011001111011101100001010000;
		#400 //2.979912e+37 * 5.576536e+20 = 5.343661e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001111101100100110000000001000;
		b = 32'b00101110000110010111111010100011;
		correct = 32'b10100001000101001011111101111001;
		#400 //-1.7589145e-29 * 3.490065e-11 = -5.039776e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011101110000110100000000001111;
		b = 32'b11001011001001010100010100001011;
		correct = 32'b00010010000101110011100000111100;
		#400 //-5.1682305e-21 * -10831115.0 = 4.7716513e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111101101001000011001001101001;
		b = 32'b00010000001100010100001000100100;
		correct = 32'b11101100111011010010001011101011;
		#400 //-0.080174275 * 3.4958048e-29 = -2.2934425e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110101001101000000000001001;
		b = 32'b00010101111111000100101010111000;
		correct = 32'b11100000001010001111001010000100;
		#400 //-4.9620908e-06 * 1.01899875e-25 = -4.869575e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100110110001001111110011000100;
		b = 32'b01110111010110011110101000101111;
		correct = 32'b10101110111001110110101001000011;
		#400 //-4.6512327e+23 * 4.4198368e+33 = -1.052354e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001100111010011001100000011001;
		b = 32'b11011111011100110011100111100100;
		correct = 32'b00101100111101011101110010110101;
		#400 //-122470600.0 * -1.752629e+19 = 6.987822e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101101111101010110110111110101;
		b = 32'b10011100100101010100010111011011;
		correct = 32'b11010000110100100111010000010000;
		#400 //2.7902106e-11 * -9.87805e-22 = -28246573000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010110010100101001100110010100;
		b = 32'b10000000001010010011100001011100;
		correct = 32'b01010110001000110111111000100110;
		#400 //-1.7012126e-25 * -3.785473e-39 = 44940550000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101111001011011001001010010101;
		b = 32'b11101101110111110011001111100101;
		correct = 32'b11000000110001110001001111000111;
		#400 //5.3718114e+28 * -8.634737e+27 = -6.221164
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011100011111100010011100010101;
		b = 32'b00000111001111000101010100001000;
		correct = 32'b11010100101011001011110000100100;
		#400 //-8.4092063e-22 * 1.4168536e-34 = -5935127000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111001100111011011001100010010;
		b = 32'b11111011000010100101011100101101;
		correct = 32'b10111110000100011110100101110101;
		#400 //1.0235282e+35 * -7.183051e+35 = -0.14249213
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100010111010100000000010110001;
		b = 32'b10001101100011101001111000110000;
		correct = 32'b11010100110100100000010010100011;
		#400 //6.342656e-18 * -8.789508e-31 = -7216167400000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100001000111000011010000001101;
		b = 32'b11001101111000011011100000000100;
		correct = 32'b01010010101100010010100010100000;
		#400 //-1.8009017e+20 * -473366660.0 = 380445400000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010111001111101010011110000101;
		b = 32'b01010001010011101011011010011000;
		correct = 32'b00000101011011000001110010111000;
		#400 //6.160375e-25 * 55489167000.0 = 1.11019415e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010101101011010111000111101;
		b = 32'b01110101100111010111011000000001;
		correct = 32'b10000100100100111011000000101100;
		#400 //-0.0013861131 * 3.9921094e+32 = -3.4721322e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001111111111001011100010111101;
		b = 32'b11000111011101111011101110010010;
		correct = 32'b00001000000000101001001111100101;
		#400 //-2.4920277e-29 * -63419.57 = 3.92943e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011110011001100011110011100010;
		b = 32'b11001000001001011100111010100001;
		correct = 32'b10010101101100011011110101000001;
		#400 //1.2188689e-20 * -169786.52 = -7.178832e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001010101101001110101101100001;
		b = 32'b01101100000001100111111111000110;
		correct = 32'b00011110001011000010110101100001;
		#400 //5928368.5 * 6.503978e+26 = 9.114988e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000111010000010111111110010101;
		b = 32'b10101001000000101101010001000110;
		correct = 32'b10011101101111010101000001011111;
		#400 //1.4557199e-34 * -2.9049916e-14 = -5.0110985e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111100111011111110110100011001;
		b = 32'b11010101011000100001001011110010;
		correct = 32'b01100111000001111101011111001000;
		#400 //-9.966143e+36 * -15535687000000.0 = 6.4149994e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110100000000011101010010010100;
		b = 32'b01111001101101010101010101100011;
		correct = 32'b00111001101101110100101000101101;
		#400 //4.114489e+31 * 1.176922e+35 = 0.00034959745
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101110011001100101101011101011;
		b = 32'b11101100100111010101100110010101;
		correct = 32'b10000001001110110110001101001000;
		#400 //5.2376697e-11 * -1.5217951e+27 = -3.4417706e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111101111100110111110011000001;
		b = 32'b10001100010010100010100100011000;
		correct = 32'b01110001000110100010101010011111;
		#400 //-0.11889029 * -1.557388e-31 = 7.633955e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110100011101011110110010011101;
		b = 32'b00001001111010001111101111001101;
		correct = 32'b01101010000001110001110000001011;
		#400 //2.2903482e-07 * 5.608876e-33 = 4.0834354e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001111100000110111001011010110;
		b = 32'b01101110001101000000101011110011;
		correct = 32'b00100000101110101110011110011001;
		#400 //4410682400.0 * 1.3930135e+28 = 3.1662884e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110001011001100110010010010000;
		b = 32'b00001010110001011001010110110100;
		correct = 32'b11100110000101010100000011111010;
		#400 //-3.3526568e-09 * 1.9026722e-32 = -1.762078e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011101011111000100111010001110;
		b = 32'b01101001111101111111111011101110;
		correct = 32'b00110011000000100011100110011111;
		#400 //1.13628905e+18 * 3.7476069e+25 = 3.032039e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100010111100111001010101001100;
		b = 32'b01010110110000101011110010001101;
		correct = 32'b10001011101000000001101101011001;
		#400 //-6.6023356e-18 * 107057540000000.0 = -6.1670906e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001000101101010111100111101111;
		b = 32'b00010111011001100001010100101111;
		correct = 32'b11110000110010011110101100011010;
		#400 //-371663.47 * 7.4343746e-25 = -4.9992566e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011010001101010110101011111010;
		b = 32'b00110010011101001001001000001101;
		correct = 32'b10100111001111011110010101100100;
		#400 //-3.7516338e-23 * 1.4235877e-08 = -2.6353372e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110110011110011100101011000010;
		b = 32'b01001101011100000001000000101000;
		correct = 32'b01101000100001010010111111111001;
		#400 //1.266596e+33 * 251724420.0 = 5.0316775e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011011110001011010101011000000;
		b = 32'b01001101001100011000101110111001;
		correct = 32'b01001110000011101000000110010110;
		#400 //1.1127662e+17 * 186170260.0 = 597714300.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010100001001001011100100101001;
		b = 32'b00010111000110001001010111111010;
		correct = 32'b01111100100010100010111010001000;
		#400 //2829924400000.0 * 4.9303146e-25 = 5.739846e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100000001000101010011001111;
		b = 32'b01111101000001011110100110100000;
		correct = 32'b00000110011111001111101000011101;
		#400 //529.32513 * 1.1125023e+37 = 4.7579686e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100000101101111010100110100011;
		b = 32'b11011101010111011000100011100100;
		correct = 32'b10000010110101000011110001101000;
		#400 //3.1113662e-19 * -9.977037e+17 = -3.1185272e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101000111000100100110001011010;
		b = 32'b00110111110110000110000001011000;
		correct = 32'b10110000100001011101111010010010;
		#400 //-2.5124153e-14 * 2.579407e-05 = -9.740282e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000011101000000000000101010001;
		b = 32'b11110001000101001101000010111111;
		correct = 32'b00010010000010011001111111100100;
		#400 //-320.01028 * -7.3689824e+29 = 4.342666e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100111110110110000111101001011;
		b = 32'b10101010010001000011001001110100;
		correct = 32'b11111101000011101110101001101100;
		#400 //2.0689607e+24 * -1.7425801e-13 = -1.1872973e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011110011101011001101010011111;
		b = 32'b00010001011101010000110000110110;
		correct = 32'b11001100100000000100101001100011;
		#400 //-1.3002167e-20 * 1.9330855e-28 = -67261210.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110100011010010001000110000111;
		b = 32'b00001000110111100100010101100111;
		correct = 32'b11101011000001100011011111001001;
		#400 //-2.1706192e-07 * 1.3377455e-33 = -1.622595e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111000111010100011110111001;
		b = 32'b10011000010101001010110001100100;
		correct = 32'b01011110001111010101001001100101;
		#400 //-9.3746285e-06 * -2.7487393e-24 = 3.4105193e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111001010001110001111001110110;
		b = 32'b00110100111111110001100111000001;
		correct = 32'b01000011110001111101001000101110;
		#400 //0.00018989466 * 4.751619e-07 = 399.64203
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001011000001110101100001100100;
		b = 32'b00100001100100111101100111111100;
		correct = 32'b10101000111010100101100010001100;
		#400 //-2.6066552e-32 * 1.0018807e-18 = -2.601762e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011010100100110110101101001110;
		b = 32'b00100111101000001100100110000110;
		correct = 32'b10110010011010101011011101000010;
		#400 //-6.0971135e-23 * 4.4627413e-15 = -1.3662261e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101100110110110100011000001000;
		b = 32'b11011010010101100010001110001111;
		correct = 32'b01010010000000110001000110110111;
		#400 //-2.1206837e+27 * -1.5068686e+16 = 140734480000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101111101001110001100101111001;
		b = 32'b00110010100100110001111111001010;
		correct = 32'b10111100100100010110000011111001;
		#400 //-3.0395222e-10 * 1.7127508e-08 = -0.017746435
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110111100000100101110111100010;
		b = 32'b01100001011011111110010000010100;
		correct = 32'b00010101100010110001111011111110;
		#400 //1.5540925e-05 * 2.7657541e+20 = 5.619055e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000010001100110111100100001000;
		b = 32'b11010111111110010110101101101101;
		correct = 32'b10101001101110000011010100110000;
		#400 //44.868195 * -548479570000000.0 = -8.180468e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001000100100000110101101100010;
		b = 32'b00001010001011110110111001011000;
		correct = 32'b11111101110100101011111011111000;
		#400 //-295771.06 * 8.446697e-33 = -3.501618e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000111001011110000010110001000;
		b = 32'b10100101110001001100111111000010;
		correct = 32'b01100000111000111010100000110010;
		#400 //-44805.53 * -3.4141362e-16 = 1.3123533e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110010011100000100110100001011;
		b = 32'b11000000010100111000101000110111;
		correct = 32'b01110001100100010110011100100110;
		#400 //-4.7596507e+30 * -3.305311 = 1.4400008e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000110101100100000101110000111;
		b = 32'b10101010101110100110100011000101;
		correct = 32'b00011011011101001000001101100010;
		#400 //-6.6973096e-35 * -3.3112936e-13 = 2.0225659e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111111001010011001011001100111;
		b = 32'b01010010011100110101011010001111;
		correct = 32'b11101100001100100110100101101111;
		#400 //-2.2542046e+38 * 261282320000.0 = -8.627468e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101010000111011100011000110110;
		b = 32'b11011101001101110000111100100111;
		correct = 32'b00001100010111001010001111100010;
		#400 //-1.401317e-13 * -8.244253e+17 = 1.69975e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111001000100111011111010111110;
		b = 32'b00111101001000101011111001101111;
		correct = 32'b01111011011010000110100000010011;
		#400 //4.794602e+34 * 0.039732393 = 1.20672375e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100100100001011011110101111100;
		b = 32'b10000000110011000100101110001100;
		correct = 32'b11100011001001111001011010100000;
		#400 //5.8000555e-17 * -1.8761542e-38 = -3.09146e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110100100001001110010100000011;
		b = 32'b00011101000011001101101001111101;
		correct = 32'b01010110111100011000100011100111;
		#400 //2.4753544e-07 * 1.8641802e-21 = 132785150000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100101001011110110101101110111;
		b = 32'b00011100010001001110111010110111;
		correct = 32'b11001000011001000000100011101011;
		#400 //-1.5215241e-16 * 6.515949e-22 = -233507.67
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011000001100110001011100101011;
		b = 32'b00000110001011110110001010111001;
		correct = 32'b11010001100000101011010000110010;
		#400 //-2.3146905e-24 * 3.2986372e-35 = -70171116000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111101001000000011011110001010;
		b = 32'b01000101000001000011110010100000;
		correct = 32'b00110111100110110001010101101011;
		#400 //0.039115466 * 2115.789 = 1.8487413e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100101010010001110101011110100;
		b = 32'b01000011111100001011101101000100;
		correct = 32'b11100000110101011010100100111100;
		#400 //-5.9300464e+22 * 481.463 = -1.2316722e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010100010010011111100110010101;
		b = 32'b01101001101100010101000011110011;
		correct = 32'b10101010000100011100110011101101;
		#400 //-3469903000000.0 * 2.6795268e+25 = -1.2949685e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011001010010101101010101010000;
		b = 32'b00010101111010000011000110011010;
		correct = 32'b11000010110111111010000100010110;
		#400 //-1.0486233e-23 * 9.378231e-26 = -111.81462
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100111111001111010111010001100;
		b = 32'b10111111001001100000011100101011;
		correct = 32'b01101000001100101001110110111001;
		#400 //-2.188173e+24 * -0.6485469 = 3.3739628e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011011010100101100011101111101;
		b = 32'b01001101101101010100000111110001;
		correct = 32'b01001101000101001101100011111000;
		#400 //5.9329085e+16 * 380124700.0 = 156077950.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010010101110101001101001111010;
		b = 32'b00110011000101000000001001111001;
		correct = 32'b00011111001000010110000001010000;
		#400 //1.1776332e-27 * 3.4461184e-08 = 3.4172744e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011100100110011100001001011011;
		b = 32'b10110110101000111111000011110100;
		correct = 32'b10100101011100000001100110110101;
		#400 //1.017493e-21 * -4.885829e-06 = -2.0825392e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001010010001100011011111110000;
		b = 32'b11101000100100001111011111010010;
		correct = 32'b00100001001011110000010010000101;
		#400 //-3247612.0 * -5.476738e+24 = 5.929829e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010000101011000110010000000110;
		b = 32'b11010111011001110110000111100011;
		correct = 32'b00111000101111101011101101100101;
		#400 //-23137890000.0 * -254407600000000.0 = 9.094811e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010011011010100001111100110100;
		b = 32'b01111001010110010011100110011111;
		correct = 32'b00011001100010011111010011011010;
		#400 //1005545850000.0 * 7.049357e+34 = 1.4264363e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111000100001100101101100010010;
		b = 32'b11110001011000001001000110001110;
		correct = 32'b00000110100110010010100100100001;
		#400 //-6.406581e-05 * -1.1120097e+30 = 5.7612637e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011001111011111001110001001;
		b = 32'b10111010001110110010011011010110;
		correct = 32'b01010000100000011110101000101101;
		#400 //-12448649.0 * -0.0007139271 = 17436862000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001111001101000110001000010011;
		b = 32'b10110001111001100110111000000001;
		correct = 32'b01011100110010000110011001011100;
		#400 //-3026326300.0 * -6.706387e-09 = 4.5126033e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111101100010010101010011111;
		b = 32'b11100110100011111100111000001101;
		correct = 32'b00010000100111011011000111101011;
		#400 //-2.1119891e-05 * -3.395497e+23 = 6.219971e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011011011011010000011000100100;
		b = 32'b10011110110000100011101010001010;
		correct = 32'b01111100000111000011001111101110;
		#400 //-6.671632e+16 * -2.056476e-20 = 3.2442063e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101111100110010011110001010110;
		b = 32'b10011000010000011101000111011100;
		correct = 32'b01010110110010100110010101011101;
		#400 //-2.787341e-10 * -2.5050617e-24 = 111268350000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010100001111011001011111110111;
		b = 32'b10101111001101110111001000111100;
		correct = 32'b01100100100001000100101000010011;
		#400 //-3257193500000.0 * -1.6684337e-10 = 1.9522463e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000001010010001011010000101001;
		b = 32'b11001110111110100110010010010010;
		correct = 32'b10110001110011010011001010111101;
		#400 //12.543984 * -2100447500.0 = -5.9720535e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100101010110011010000101011001;
		b = 32'b01011000010011000111111101111100;
		correct = 32'b00001100100010000011100001000101;
		#400 //1.8876416e-16 * 899391650000000.0 = 2.0987984e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110111001111011111000111001100;
		b = 32'b01111111011110011010110001111100;
		correct = 32'b10110111010000101100000111100001;
		#400 //-3.8525325e+33 * 3.3187336e+38 = -1.1608442e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001110110100111011111100101110;
		b = 32'b00001000101000100100111100111000;
		correct = 32'b01000101101001101111110010110101;
		#400 //5.2199615e-30 * 9.768645e-34 = 5343.5884
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000000010110110010101000000010;
		b = 32'b00101110101111100001110010101111;
		correct = 32'b00010000111101011000010010111001;
		#400 //8.3721e-39 * 8.645295e-11 = 9.683995e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011011001011010010000111101110;
		b = 32'b10110101010100000000010011011011;
		correct = 32'b11100101010101010001000100011000;
		#400 //4.8732477e+16 * -7.7493104e-07 = -6.288621e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001000001101000111010101001010;
		b = 32'b01000000011011001000100010011010;
		correct = 32'b00000111010000110100111101000100;
		#400 //5.4304652e-34 * 3.6958375 = 1.4693464e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110010011111011111001101110101;
		b = 32'b01100100010111001110110100011000;
		correct = 32'b10001101100100110010001001001000;
		#400 //-1.4781894e-08 * 1.6301472e+22 = -9.067827e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010000100010011111101100000100;
		b = 32'b11010111011100111000001100010010;
		correct = 32'b10111000100100010000111001111100;
		#400 //18519433000.0 * -267744270000000.0 = -6.916837e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011100100011000100110010100111;
		b = 32'b01111100010000100110101011101101;
		correct = 32'b00011111101110001011110101011001;
		#400 //3.159262e+17 * 4.0378972e+36 = 7.824028e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000101111110000000101101001011;
		b = 32'b01010010101001111010110010011011;
		correct = 32'b00110010101111010101101001101000;
		#400 //7937.4116 * 360077700000.0 = 2.2043608e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111001100000100000100101001101;
		b = 32'b00111001010110100000100110110000;
		correct = 32'b00111111100110001010110100111101;
		#400 //0.00024802462 * 0.00020793709 = 1.1927868
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110011110111001101011111001111;
		b = 32'b00010100110100100101001010010010;
		correct = 32'b11011110100001100110011100010011;
		#400 //-1.0283804e-07 * 2.123715e-26 = -4.842365e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011101001100110100111101011011;
		b = 32'b10011011011111110001100010001101;
		correct = 32'b11000001001100111111001000001011;
		#400 //2.3731479e-21 * -2.1101038e-22 = -11.2465925
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101001001101111111111100000110;
		b = 32'b00110110010100111011000101000110;
		correct = 32'b11110010010111101000000111000000;
		#400 //-1.3902359e+25 * 3.1544637e-06 = -4.407202e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000011011100000011111001010000;
		b = 32'b10011010111101101110000001110011;
		correct = 32'b01100111111110010001111100011100;
		#400 //-240.24341 * -1.0210583e-22 = 2.3528862e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100011110101001110001100010000;
		b = 32'b11000111100111110110101100000001;
		correct = 32'b01011011101010101110111001101101;
		#400 //-7.8541426e+21 * -81622.01 = 9.62258e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101110100010111010000000010111;
		b = 32'b00111100011001111000000101100110;
		correct = 32'b10110001100110100110011000000010;
		#400 //-6.349426e-11 * 0.014129972 = -4.493587e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110110110010110111001101000101;
		b = 32'b01001101011101100100110001010100;
		correct = 32'b00101000110100110111011011011101;
		#400 //6.0632906e-06 * 258262340.0 = 2.3477255e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001011110110110001000000110010;
		b = 32'b11000011100000001011110010011001;
		correct = 32'b11000111110110011100111101000101;
		#400 //28713060.0 * -257.47342 = -111518.54
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110110101111000000101001111;
		b = 32'b11100111111000111000010110011101;
		correct = 32'b10010110011100100111101010100101;
		#400 //0.42090842 * -2.1488838e+24 = -1.9587304e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100000000101111100011101100001;
		b = 32'b11000101111110010110110000111111;
		correct = 32'b00011001100110111100011111111010;
		#400 //-1.2856166e-19 * -7981.531 = 1.6107394e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111111110010110011101111001010;
		b = 32'b01100000110010000011010111001011;
		correct = 32'b00011110100000011110111011010110;
		#400 //1.5877621 * 1.1541328e+20 = 1.3757187e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111000011001000100010001011011;
		b = 32'b00101011100100001101000001100111;
		correct = 32'b01001100010010011100001101101101;
		#400 //5.4423097e-05 * 1.0289659e-12 = 52891060.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001001011110000111010000001011;
		b = 32'b00000110001001010110011101011000;
		correct = 32'b01000010110000000100010011100101;
		#400 //2.9906477e-33 * 3.1108976e-35 = 96.13456
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111111100110100111111001111101;
		b = 32'b11111100110000001001001110111110;
		correct = 32'b00000010010011010101111111110011;
		#400 //-1.2069851 * -7.9993405e+36 = 1.5088557e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111000001000110110111001001110;
		b = 32'b00011100010101110011000001011111;
		correct = 32'b11011011010000100110110100001000;
		#400 //-3.8964958e-05 * 7.120005e-22 = -5.4726027e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001001101010100011001010010111;
		b = 32'b10100100010101110011100100001010;
		correct = 32'b11100100110010100111000110110001;
		#400 //1394258.9 * -4.6669007e-17 = -2.9875477e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101111101001010111001110010010;
		b = 32'b00100110000010010100010110110011;
		correct = 32'b11001001000110100100011010011001;
		#400 //-3.0095443e-10 * 4.7625883e-16 = -631913.56
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001101001101001001011111101000;
		b = 32'b00100111001111110100111010110110;
		correct = 32'b01100101011100011010100110110000;
		#400 //189365890.0 * 2.6549244e-15 = 7.132628e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011010111011001101100110010101;
		b = 32'b11001011100010110110010101001010;
		correct = 32'b00001110110110010111110011000010;
		#400 //-9.7958835e-23 * -18270868.0 = 5.3614768e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111000100100101001101111001001;
		b = 32'b10100000101001000111110110111100;
		correct = 32'b11010111011001000010101101000101;
		#400 //6.99084e-05 * -2.7865885e-19 = -250874500000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110100001011010010110100001000;
		b = 32'b11100111011001000010101101001110;
		correct = 32'b01001100010000100100110010001001;
		#400 //-5.4881634e+31 * -1.0774984e+24 = 50934308.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001110010011010001011111100001;
		b = 32'b10001011101110100101111001100110;
		correct = 32'b01000010000011001101110000110110;
		#400 //-2.5279698e-30 * -7.178663e-32 = 35.21505
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000011011000110101111101100010;
		b = 32'b00010001101110100111010111100110;
		correct = 32'b00110001000111000001010111000010;
		#400 //6.68188e-37 * 2.9418286e-28 = 2.2713356e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111011001110011100010110100010;
		b = 32'b10100010011010000100100001111110;
		correct = 32'b11011000010011001011110101101010;
		#400 //0.0028346558 * -3.148024e-18 = -900455600000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000111100111111100111110011010;
		b = 32'b10111111010011101101111101100011;
		correct = 32'b10000111110001011100001100100110;
		#400 //2.4045678e-34 * -0.8080961 = -2.9755963e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010011010111111010101110100011;
		b = 32'b00000101000101000000010101111010;
		correct = 32'b01001101110000010110101010110001;
		#400 //2.823118e-27 * 6.9599324e-36 = 405624350.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000011010111110010000001000111;
		b = 32'b10011001101000010000111111100001;
		correct = 32'b10101001001100010101001011101000;
		#400 //6.5570863e-37 * -1.6653423e-23 = -3.9373805e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111111101101010100010100110000;
		b = 32'b10101000110111000010101001010001;
		correct = 32'b01010110010100101100011000111001;
		#400 //-1.4161739 * -2.4443258e-14 = 57937200000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010111010101000110100100110;
		b = 32'b01000110110000010011110010100100;
		correct = 32'b10110011100110110101110111011111;
		#400 //-0.0017894849 * 24734.32 = -7.234825e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111001010010101111101100010010;
		b = 32'b11001000001100010100100101111011;
		correct = 32'b00110000100100101000110011111001;
		#400 //-0.00019357752 * -181541.92 = 1.0662965e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010101011000101000010111110;
		b = 32'b11110111011100111010001000101001;
		correct = 32'b00000010101101010000111111011011;
		#400 //-0.0013146622 * -4.9414732e+33 = 2.660466e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111010110001001110101010111001;
		b = 32'b01000110010111001111001010100101;
		correct = 32'b00110011111001000010100000011100;
		#400 //0.0015023566 * 14140.661 = 1.0624373e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110110001110011100101001010110;
		b = 32'b11010010101110111100100001001010;
		correct = 32'b10100010111111010100100011001010;
		#400 //2.7684923e-06 * -403259600000.0 = -6.8652856e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000011000100111110010000101011;
		b = 32'b10100010110100101100111100010111;
		correct = 32'b11011111101100111001100000111110;
		#400 //147.89128 * -5.713988e-18 = -2.5882323e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001100010010111010100000000011;
		b = 32'b10011111100000110110111110101111;
		correct = 32'b01101100010001100101010011111000;
		#400 //-53387276.0 * -5.566542e-20 = 9.590743e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001000010101000110000001011110;
		b = 32'b00010100100010010111010110111001;
		correct = 32'b11110011010001011100001011001010;
		#400 //-217473.47 * 1.3879898e-26 = -1.5668232e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100111110010011111010110111111;
		b = 32'b00110100001011010101010101011101;
		correct = 32'b10110011000101010010001110111010;
		#400 //-5.6055145e-15 * 1.6142936e-07 = -3.472426e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100100100111101100100000000110;
		b = 32'b00101111111010010001010111100001;
		correct = 32'b11110100001011100110010000011101;
		#400 //-2.343199e+22 * 4.2398e-10 = -5.5266735e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111111010001111000001000100110;
		b = 32'b00111001101001000110000101000100;
		correct = 32'b11000101000110110101101010011101;
		#400 //-0.77932966 * 0.00031352986 = -2485.6633
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100100011011110111010111001010;
		b = 32'b00010101000111011010011101111010;
		correct = 32'b01001110110000100110101100100011;
		#400 //5.1924635e-17 * 3.1838013e-26 = 1630900600.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010110010001011101111010100111;
		b = 32'b10101000100010010111111100000010;
		correct = 32'b10101101001110000011010000110101;
		#400 //1.598379e-25 * -1.5265136e-14 = -1.0470781e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001001000000111100000111011010;
		b = 32'b01111110110111111110000110110101;
		correct = 32'b10001001100101101010100011000111;
		#400 //-539677.6 * 1.4879489e+38 = -3.6269904e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001100000101000000001110011101;
		b = 32'b10101001011011000101110011111010;
		correct = 32'b11100010001000000100111110011100;
		#400 //38801012.0 * -5.248317e-14 = -7.393039e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111001100010000010110111111010;
		b = 32'b01101010011001101110000011001100;
		correct = 32'b01001110100101101111111101010000;
		#400 //8.838561e+34 * 6.977863e+25 = 1266657300.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000100000101000010001000101111;
		b = 32'b01001110011101010100101010100110;
		correct = 32'b10110101000110101001100110110101;
		#400 //-592.5341 * 1028827500.0 = -5.7593144e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100100000101000000000101000011;
		b = 32'b10101101100111110001100011111100;
		correct = 32'b01110101111011100010011010101100;
		#400 //-1.0920836e+22 * -1.8087302e-11 = 6.0378467e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111010010100000011100000110011;
		b = 32'b11010111100000111111010101001110;
		correct = 32'b01100010010010011111100101001001;
		#400 //-2.702844e+35 * -290179200000000.0 = 9.314396e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111000110001101100100001100110;
		b = 32'b10011001110010011011001010111011;
		correct = 32'b11011110011111000100110010111101;
		#400 //9.478703e-05 * -2.0855102e-23 = -4.5450284e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010110010011100110010101010111;
		b = 32'b11110011001000011110010100110110;
		correct = 32'b10100010101000110010111100000010;
		#400 //56733660000000.0 * -1.2826672e+31 = -4.423101e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001001101001011100011111101001;
		b = 32'b11110111010101001010001111011010;
		correct = 32'b00010001110001111001010111110000;
		#400 //-1358077.1 * -4.3128525e+33 = 3.148907e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111011100110001000101010100011;
		b = 32'b00111010001010011110111010001111;
		correct = 32'b01000000111001011100110100111110;
		#400 //0.0046551987 * 0.00064823864 = 7.181304
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100100101111011011001011001001;
		b = 32'b11001100000101000000111100100110;
		correct = 32'b01011000001000111111111101110110;
		#400 //-2.799454e+22 * -38812824.0 = 721270400000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111001101011011111100010101011;
		b = 32'b11000000010010110010111000100111;
		correct = 32'b11111000110110110011001010100010;
		#400 //1.1291387e+35 * -3.174692 = -3.5566874e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100111011010011011101010110001;
		b = 32'b10001100000010011100101110101100;
		correct = 32'b01011010110110010001110100101100;
		#400 //-3.2436451e-15 * -1.0615386e-31 = 3.0556072e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101100000110100101011111011001;
		b = 32'b01101000101100001111100101000000;
		correct = 32'b00000010110111110100001110011000;
		#400 //2.1933482e-12 * 6.685875e+24 = 3.2805702e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100001011110011001010111100110;
		b = 32'b00001101101110011000010011010011;
		correct = 32'b01010011001011000011010000001001;
		#400 //8.456287e-19 * 1.1433482e-30 = 739607400000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010001100111001100000101110000;
		b = 32'b01010000111011010000011000010101;
		correct = 32'b01000000001010010100111000111000;
		#400 //84157530000.0 * 31812790000.0 = 2.645399
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101101011100111100010001111001;
		b = 32'b10010000011011111010011101000010;
		correct = 32'b01011100100000100011001010000111;
		#400 //-1.38565765e-11 * -4.726329e-29 = 2.9317842e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010001000110101010100111000000;
		b = 32'b00111111000011000110110110100100;
		correct = 32'b00010001100011001111100110011001;
		#400 //1.2200766e-28 * 0.548548 = 2.2241932e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111001111110101100001010000110;
		b = 32'b11110100010110011100001001101101;
		correct = 32'b01000101000100110110010111010100;
		#400 //-1.6275245e+35 * -6.9010733e+31 = 2358.3643
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110110000011101010010111101100;
		b = 32'b11100110100110111100101110010100;
		correct = 32'b01001110111010100110010110011101;
		#400 //-7.23312e+32 * -3.6786108e+23 = 1966263900.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001110101101000010101100001100;
		b = 32'b01101011100010000100101010101111;
		correct = 32'b10100010101010010011010100000010;
		#400 //-1511360000.0 * 3.295332e+26 = -4.5863666e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001010011000101111000011011111;
		b = 32'b11100111111010100100101100001001;
		correct = 32'b10100001111101111111011101110101;
		#400 //3718199.8 * -2.2128358e+24 = -1.6802872e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101111100000111110100101000110;
		b = 32'b00100001011011100011011110111000;
		correct = 32'b01001101100011011100001000010001;
		#400 //2.3994512e-10 * 8.071128e-19 = 297288220.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010101010111101011011111110;
		b = 32'b01101110101011110001010011000101;
		correct = 32'b10001011011110110100001010110111;
		#400 //-0.0013110337 * 2.7092493e+28 = -4.8391032e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110101100100101100011010100101;
		b = 32'b01011100001111000000010010100011;
		correct = 32'b10011000110001111101100010001011;
		#400 //-1.0935661e-06 * 2.1168957e+17 = -5.1658947e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011001010000100000111101011101;
		b = 32'b11110110110101011111011001011100;
		correct = 32'b10100001111010000010111111111011;
		#400 //3413939800000000.0 * -2.169836e+33 = -1.5733632e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001011001111110010011100011110;
		b = 32'b01110101001000111111100010111001;
		correct = 32'b00010101100101010011011111100010;
		#400 //12527390.0 * 2.0785866e+32 = 6.026879e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100110101000010000001000010;
		b = 32'b01001111000000000010001110000110;
		correct = 32'b00110101010100111110010101110011;
		#400 //1697.008 * 2149811700.0 = 7.893752e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101000100001100111011011000011;
		b = 32'b11101010101101100010111001101011;
		correct = 32'b10111101001111001111001010100100;
		#400 //5.079903e+24 * -1.1012185e+26 = -0.046129838
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011001100011100000001110001011;
		b = 32'b11001010001011101000011000000000;
		correct = 32'b00001110110100000101000000110001;
		#400 //-1.4683887e-23 * -2859392.0 = 5.135318e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000001010100001011001000011;
		b = 32'b11101010100110011011111101011000;
		correct = 32'b00000101000011011001101001101100;
		#400 //-6.1877276e-10 * -9.293462e+25 = 6.658151e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101001001111011100000000010100;
		b = 32'b00010100010010101110000001100101;
		correct = 32'b01010100011011110110111111001000;
		#400 //4.213303e-14 * 1.0242648e-26 = 4113490200000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111110001110000101011001100000;
		b = 32'b11011000001110001100100100000011;
		correct = 32'b00100101011111110110000100101111;
		#400 //-0.180017 * -812693900000000.0 = 2.2150651e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110100011000010001101111100011;
		b = 32'b11111111111011110011001110000111;
		correct = 32'b11111111111011110011001110000111;
		#400 //-7.133987e+31 * nan = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001010101000100011110110101001;
		b = 32'b00110000101001010101000000110011;
		correct = 32'b10011001011110110011110111111100;
		#400 //-1.5623227e-32 * 1.2028124e-09 = -1.29889135e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100101101100111101010011101010;
		b = 32'b10010000000000101100010000110000;
		correct = 32'b01010101001100000000011100000001;
		#400 //-3.1195826e-16 * -2.5789117e-29 = 12096508000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011110010110101110010011000001;
		b = 32'b10110000000000100000011001110001;
		correct = 32'b01101101110101110111101111111001;
		#400 //-3.943236e+18 * -4.730288e-10 = 8.336144e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011010110110011110011101000100;
		b = 32'b11010011001111110110011100001010;
		correct = 32'b10000111000100011011100011110000;
		#400 //9.0122726e-23 * -822067460000.0 = -1.0962936e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110011111111110011001001100110;
		b = 32'b00111001001000110110111100100000;
		correct = 32'b11111010010001111101111000100100;
		#400 //-4.0437558e+31 * 0.00015586289 = -2.5944316e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101111111101001111110101101110;
		b = 32'b11001001011100001010100001001110;
		correct = 32'b00100110000000100100110111101011;
		#400 //-4.4563414e-10 * -985732.9 = 4.520841e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001011101100000101010110110001;
		b = 32'b00010010000111111100000111000110;
		correct = 32'b01111001000011010100100001001101;
		#400 //23112546.0 * 5.04104e-28 = 4.584877e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000000000011111111011100111101;
		b = 32'b00011111101001011110010010001001;
		correct = 32'b01011111110111100010100111000000;
		#400 //2.2494652 * 7.02583e-20 = 3.2017075e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000100000110101100010100010000;
		b = 32'b10011100101101100011011000000001;
		correct = 32'b10100110110110010111001000110100;
		#400 //1.81931e-36 * -1.2057709e-21 = -1.5088355e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101011011111000000001010111100;
		b = 32'b10101011000001011110101010101001;
		correct = 32'b00111111111100001110000001100000;
		#400 //-8.953218e-13 * -4.757675e-13 = 1.8818474
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110010111010110110011001000;
		b = 32'b01011110101001011111010001000101;
		correct = 32'b10010111001010101100100011010001;
		#400 //-3.2994885e-06 * 5.9791294e+18 = -5.518343e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110111010111100100101000110000;
		b = 32'b01100010000000110010000100100100;
		correct = 32'b11010100110110001111110000011001;
		#400 //-4.5085727e+33 * 6.047279e+20 = -7455539500000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001010111111011000111110010110;
		b = 32'b10101100111101001110000100101010;
		correct = 32'b10011101100001001000100110101100;
		#400 //2.4417025e-32 * -6.9598953e-12 = -3.508246e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100000100110010101011010011110;
		b = 32'b00100100011000110001010110010111;
		correct = 32'b00111011101011001101110100010101;
		#400 //2.5976527e-19 * 4.9241066e-17 = 0.0052753785
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110011010110110110001100101000;
		b = 32'b11001010111010100001100110111000;
		correct = 32'b11100111111011111110100100010110;
		#400 //1.7381655e+31 * -7671004.0 = -2.2658905e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100001000101110110000111111010;
		b = 32'b01001101110110001000111001100010;
		correct = 32'b00010010101100101111010010101101;
		#400 //5.129046e-19 * 454151230.0 = 1.1293697e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000110000110101110001111001000;
		b = 32'b10100101001011000100010110100000;
		correct = 32'b01100000011001100010101101101111;
		#400 //-9912.945 * -1.4942212e-16 = 6.634189e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100100000010000110001110010010;
		b = 32'b10101011011100100100010101001010;
		correct = 32'b00111000000100000001111000110111;
		#400 //-2.957464e-17 * -8.607183e-13 = 3.4360415e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000100011001110000000010000010;
		b = 32'b00101110111001011100000000000011;
		correct = 32'b10010101000000001011001010001111;
		#400 //-2.7154153e-36 * 1.04478225e-10 = -2.5990252e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101010111101101111100000001100;
		b = 32'b11110100111011010100011000100011;
		correct = 32'b10110101100001010011101011100101;
		#400 //1.4928356e+26 * -1.5039025e+32 = -9.926413e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110111110111001100100110011110;
		b = 32'b01111011111000111111110010001011;
		correct = 32'b10111011011101111110101010100001;
		#400 //-8.956208e+33 * 2.3675471e+36 = -0.0037829059
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011101011000100111100001010101;
		b = 32'b00111111000101011111101000001111;
		correct = 32'b10011101110000010100100011001011;
		#400 //-2.9973061e-21 * 0.58584684 = -5.116194e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000110111100110001111000010000;
		b = 32'b00110000111101100100001011101100;
		correct = 32'b01010101011111001011101101010000;
		#400 //31119.031 * 1.7917876e-09 = 17367589000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110010110111111000101111001001;
		b = 32'b10101110101000100001011111111100;
		correct = 32'b01000011101100001000011011100001;
		#400 //-2.6024184e-08 * -7.3711676e-11 = 353.05374
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101101110111000101000101001101;
		b = 32'b11010000000100000100100000100001;
		correct = 32'b01011101010000110111010010010110;
		#400 //-8.5231236e+27 * -9682585000.0 = 8.802529e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111100100111100011111101111010;
		b = 32'b01010100111010111100000100110100;
		correct = 32'b00100111001010111101011001100000;
		#400 //0.019317377 * 8100470000000.0 = 2.384723e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000000010010100110100101010000;
		b = 32'b00111000101111001010011011011100;
		correct = 32'b10000110110010011111001110111100;
		#400 //-6.833606e-39 * 8.9956186e-05 = -7.596593e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010011110101001000011000001010;
		b = 32'b00011001111111001111100110100100;
		correct = 32'b10111001010101110001000010010011;
		#400 //-5.3648497e-27 * 2.6157018e-23 = -0.00020510172
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111110010111000100101001101010;
		b = 32'b11000001001110011100100100110010;
		correct = 32'b00111100100101111100010111000111;
		#400 //-0.21512762 * -11.61162 = 0.018526925
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100001010010100101100101110101;
		b = 32'b00001001000100110101000100101101;
		correct = 32'b01010111101011111101000011110001;
		#400 //6.855866e-19 * 1.773265e-33 = 386623860000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110100110111101011100011000;
		b = 32'b11011101011011101100011101111111;
		correct = 32'b10100000101001110001010001010010;
		#400 //0.3043754 * -1.0753663e+18 = -2.8304347e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110010110101110001111110101111;
		b = 32'b01101100110010101110111111110111;
		correct = 32'b11000101100001111010111110111000;
		#400 //-8.52193e+30 * 1.9626897e+27 = -4341.965
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111011110111110101101011001100;
		b = 32'b01001100000101101110001000011110;
		correct = 32'b01101111001111010111101011110001;
		#400 //2.3194476e+36 * 39553144.0 = 5.8641294e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110001111111000110110110010100;
		b = 32'b00100100001000011110011011001011;
		correct = 32'b01001101010001111001001000010100;
		#400 //7.346623e-09 * 3.51068e-17 = 209264960.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101101011000100001100001001001;
		b = 32'b11100001011101011110000111111101;
		correct = 32'b10001011011010110110010111011100;
		#400 //1.2852005e-11 * -2.8348353e+20 = -4.5335984e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111000110101000101101100001001;
		b = 32'b01011010100011011100101011001011;
		correct = 32'b11011101101111111011001100100001;
		#400 //-3.4456667e+34 * 1.9955472e+16 = -1.7266776e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110011111010100100000111100;
		b = 32'b11100100110011111101000000011001;
		correct = 32'b00010001000111000000000110011100;
		#400 //-3.7741984e-06 * -3.0667768e+22 = 1.2306726e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010000101111100000101101010011;
		b = 32'b10010101101010100011001101110111;
		correct = 32'b01111010100011101110110001010001;
		#400 //-25507305000.0 * -6.874365e-26 = 3.710496e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111110100011001000101010101111;
		b = 32'b10000011001011000001000101110110;
		correct = 32'b01111010110100010001100001110001;
		#400 //-0.27449557 * -5.05663e-37 = 5.428429e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010110011100011010011111101100;
		b = 32'b11000010111101001100100111010010;
		correct = 32'b11010010111111001011100101100000;
		#400 //66425880000000.0 * -122.39418 = -542720920000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001001001011111001001100010001;
		b = 32'b10100110100101110011110110110110;
		correct = 32'b10100010000101001001100000011001;
		#400 //2.1134009e-33 * -1.0494457e-15 = -2.013826e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000001110100101000001001101010;
		b = 32'b10110111100100101001100110010000;
		correct = 32'b11001001101101111100110100010010;
		#400 //26.313679 * -1.7476064e-05 = -1505698.2
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000101101111000101001100100011;
		b = 32'b00011000101000110011000111011100;
		correct = 32'b01101100100100111011010111011111;
		#400 //6026.392 * 4.2184858e-24 = 1.4285677e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011101010011011111001010000110;
		b = 32'b00010010011100100111111101000010;
		correct = 32'b01001010010110010110101001000010;
		#400 //2.7256906e-21 * 7.6518593e-28 = 3562128.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111100010010011101101010010011;
		b = 32'b11000011101011001110010101101110;
		correct = 32'b11111000000101010111000000101010;
		#400 //4.1923395e+36 * -345.79242 = -1.2123862e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110001100100111001111000101000;
		b = 32'b01001100011000110000110110001101;
		correct = 32'b10100100101001100111000000001010;
		#400 //-4.2962434e-09 * 59520564.0 = -7.2180826e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101001000010011000100001000001;
		b = 32'b11000111011001111100101011111110;
		correct = 32'b00100001000101111110010100110001;
		#400 //-3.0538292e-14 * -59338.992 = 5.146412e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100010111100101110011000100101;
		b = 32'b10100011100101010111110110010111;
		correct = 32'b00111110110011111111101011101010;
		#400 //-6.5837906e-18 * -1.6207802e-17 = 0.4062112
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000010011011111000001011011001;
		b = 32'b01100110100011000011110000000001;
		correct = 32'b00011011010110101001110110010111;
		#400 //59.87778 * 3.311191e+23 = 1.8083457e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011000010100111111000100000111;
		b = 32'b11010111000000001100111010100010;
		correct = 32'b11000000110100101001110100001000;
		#400 //932128600000000.0 * -141624970000000.0 = -6.581669
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001011001111011100001101110010;
		b = 32'b00000001100011101011000000100110;
		correct = 32'b11001001001010100011101011000010;
		#400 //-3.6547113e-32 * 5.241532e-38 = -697260.1
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111000010000110011001110101000;
		b = 32'b11100110110010111001001001110111;
		correct = 32'b11010000111101010111100101010101;
		#400 //1.583665e+34 * -4.806711e+23 = -32946956000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101111101100011000101100100011;
		b = 32'b11010011000000011100110111011010;
		correct = 32'b11011100001011110001001101101101;
		#400 //1.0989411e+29 * -557504400000.0 = -1.9711792e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111001001010010111000111010110;
		b = 32'b10010100100101000010010001010101;
		correct = 32'b01100100000100100110100000000111;
		#400 //-0.00016159503 * -1.4958511e-26 = 1.0802882e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111010010111001001011011010101;
		b = 32'b01010100111110011001000110000110;
		correct = 32'b01100100111000100100011000100000;
		#400 //2.8634114e+35 * 8575106700000.0 = 3.3392138e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100101010100110010001010000001;
		b = 32'b11111100100001110101011101000000;
		correct = 32'b10101000010001111010111011010101;
		#400 //6.231599e+22 * -5.621838e+36 = -1.108463e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110110110100000011011101111000;
		b = 32'b01000011111001010100100100110101;
		correct = 32'b01110010011010000111100111010111;
		#400 //2.111568e+33 * 458.57193 = 4.6046603e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000011100010011000111100110001;
		b = 32'b10001010111001000001100011001011;
		correct = 32'b11111000000110100110001100010011;
		#400 //275.11868 * -2.1964927e-32 = -1.2525362e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011100001101110100100101110010;
		b = 32'b00101111111111001100101111111001;
		correct = 32'b00101011101110011001101111111111;
		#400 //6.0644547e-22 * 4.5983464e-10 = 1.3188338e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011001011101000101101111011110;
		b = 32'b11010101100001101010101101111011;
		correct = 32'b11000011011010000100000110100011;
		#400 //4298806500000000.0 * -18508883000000.0 = -232.2564
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110111110010001111001100011001;
		b = 32'b11011101011111101000110000111010;
		correct = 32'b01011001110010100001100010010111;
		#400 //-8.151484e+33 * -1.1463812e+18 = 7110623000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100110111001101110011100111001;
		b = 32'b01010110011101011001011110101001;
		correct = 32'b00001111111100001011000000110100;
		#400 //1.6022129e-15 * 67507930000000.0 = 2.3733698e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110100111001010011111010011110;
		b = 32'b01101110101101001010110001101010;
		correct = 32'b01000101101000100110100100100100;
		#400 //1.4530103e+32 * 2.7957869e+28 = 5197.1426
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011100000110100011001001101010;
		b = 32'b10101101011011001101101101100111;
		correct = 32'b01101110001001101010100011000100;
		#400 //-1.7361031e+17 * -1.3463764e-11 = 1.2894634e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011100001111001001110100100001;
		b = 32'b01000011010101101010000010100000;
		correct = 32'b11011000011000001111100011001010;
		#400 //-2.1236024e+17 * 214.62744 = -989436600000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100110011101111001000000111111;
		b = 32'b00010000011000110111111001111010;
		correct = 32'b01010101100010110100101011000111;
		#400 //8.589083e-16 * 4.486529e-29 = 19144160000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011111100100110010110100010010;
		b = 32'b10011011000100111100100010110000;
		correct = 32'b01000011111111101111001001101110;
		#400 //-6.2331484e-20 * -1.2224401e-22 = 509.89398
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111000100100001101100111000111;
		b = 32'b11001110000010000011100001011110;
		correct = 32'b00101010000010000001110000010101;
		#400 //-6.907019e-05 * -571348860.0 = 1.208897e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100001111110001011101100110111;
		b = 32'b00000001111001100000101100001011;
		correct = 32'b01011111100010100110010111111111;
		#400 //1.6854689e-18 * 8.45045e-38 = 1.9945315e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100111010011100100101011101100;
		b = 32'b11001110111000111111110100111111;
		correct = 32'b00010111111001111010001101000110;
		#400 //-2.8628858e-15 * -1912512400.0 = 1.4969241e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101000001001000110010111101000;
		b = 32'b00101000111011111100100101011001;
		correct = 32'b10111110101011111000001110011010;
		#400 //-9.125926e-15 * 2.6621651e-14 = -0.34280092
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111111010001110010000100100111;
		b = 32'b11111000010111100101111011100110;
		correct = 32'b11000110011001010011111001111000;
		#400 //2.646885e+38 * -1.8040854e+34 = -14671.617
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110001010011100111110010000001;
		b = 32'b01101101110111100011011100000101;
		correct = 32'b01000010111011011110000101001101;
		#400 //1.02247085e+30 * 8.5965233e+27 = 118.94004
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010011010101110011110111111;
		b = 32'b01111000101011010110100000111101;
		correct = 32'b10000001001011010110010100000110;
		#400 //-0.00089609245 * 2.8136924e+34 = -3.1847562e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010100000110111000101100111110;
		b = 32'b00111010111111110111001101111010;
		correct = 32'b10011000100110111110000011001111;
		#400 //-7.852961e-27 * 0.0019489371 = -4.029356e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000000100000011000000110110010;
		b = 32'b00011001110100000100001010110010;
		correct = 32'b10100110000111110011000110000001;
		#400 //-1.1893305e-38 * 2.1533634e-23 = -5.5231297e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010011000010110100001001000001;
		b = 32'b11100110001000011011000101111100;
		correct = 32'b10101100010111000111101100010000;
		#400 //598112000000.0 * -1.9089375e+23 = -3.1332194e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100010010010101100011111010011;
		b = 32'b11011011101100110010001001110101;
		correct = 32'b01000110000100001110010101101010;
		#400 //-9.351603e+20 * -1.0084381e+17 = 9273.354
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000001101001101000001110111011;
		b = 32'b10011110100110110000100100101011;
		correct = 32'b11100010100010010111101000100000;
		#400 //20.814322 * -1.6415055e-20 = -1.268002e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101011101111010100111111010100;
		b = 32'b01101110101100011010111001001101;
		correct = 32'b10111100100010000110000011111101;
		#400 //-4.577279e+26 * 2.7494782e+28 = -0.01664781
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011101010011010101011010011111;
		b = 32'b00100000101010010110110001100011;
		correct = 32'b00111100000110110010001001000111;
		#400 //2.7176306e-21 * 2.8701438e-19 = 0.009468622
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011011010101011111111111001001;
		b = 32'b11001001010110111011110001101011;
		correct = 32'b01010001011110010101000011111110;
		#400 //-6.023541e+16 * -900038.7 = 66925355000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011000110011001000011011000100;
		b = 32'b11011100010100001001101100110110;
		correct = 32'b10111011111110101111111001000100;
		#400 //1799033500000000.0 * -2.348698e+17 = -0.0076597054
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010010110101111101000000011011;
		b = 32'b11100010101011100100000111110000;
		correct = 32'b10101111100111101000011000110110;
		#400 //463454700000.0 * -1.6072424e+21 = -2.8835395e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001000001111010001001111111101;
		b = 32'b10011001001100110101010001100110;
		correct = 32'b10101110100001101111010101000110;
		#400 //5.6898615e-34 * -9.271127e-24 = -6.137184e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100101000001010010101111010010;
		b = 32'b11111011010010100110100010101110;
		correct = 32'b10101001001010000110111000110001;
		#400 //3.9305193e+22 * -1.0509671e+36 = -3.739907e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110011111000110111010010110110;
		b = 32'b10010101100111111001010000010000;
		correct = 32'b01011101101101100111001000001100;
		#400 //-1.0591741e-07 * -6.445319e-26 = 1.643323e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101001111101111100001110100100;
		b = 32'b11011111000010010010011101111001;
		correct = 32'b01001010011001110011101000111101;
		#400 //-3.744107e+25 * -9.883001e+18 = 3788431.2
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101110110111011010100101111000;
		b = 32'b10111110100110011010010110001110;
		correct = 32'b11101111101110001010100110000101;
		#400 //3.430053e+28 * -0.3000912 = -1.1430036e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001000100100100000111111101000;
		b = 32'b00001101110111110000011011010110;
		correct = 32'b01111010001001111010100000011001;
		#400 //299135.25 * 1.3745082e-30 = 2.1763075e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010111000111000010110001100011;
		b = 32'b10100001010011011101010010000000;
		correct = 32'b11110101010000100011110101100001;
		#400 //171714450000000.0 * -6.9737943e-19 = -2.4622815e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010011111010000101011010010001;
		b = 32'b00110101100001011011011111001100;
		correct = 32'b10011101110111100110011100101111;
		#400 //-5.8650395e-27 * 9.962764e-07 = -5.88696e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010000001110111000001100110010;
		b = 32'b01101100011110101110001100011110;
		correct = 32'b10100011001111110101010101110100;
		#400 //-12583750000.0 * 1.21321594e+27 = -1.0372226e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111100100101010001111011111101;
		b = 32'b00001000101010000111000110101111;
		correct = 32'b11110011011000101010001000001101;
		#400 //-0.018203253 * 1.0137859e-33 = -1.7955717e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010111010101101011101111000001;
		b = 32'b10011001000010000100000010110110;
		correct = 32'b10111101110010011011101000100011;
		#400 //6.938411e-25 * -7.0441035e-24 = -0.09849956
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101100101110111101100100000000;
		b = 32'b11000110011000100101010011111110;
		correct = 32'b10100101110101000111100010010111;
		#400 //5.3389515e-12 * -14485.248 = -3.6857853e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011011000000110100111101111100;
		b = 32'b01111000101011110000011110011111;
		correct = 32'b00100001110000000000111001001010;
		#400 //3.6960616e+16 * 2.8400204e+34 = 1.3014208e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111011111010101100101100010111;
		b = 32'b00001011001111011000000010111001;
		correct = 32'b01110000000111101001011101101111;
		#400 //0.0071653235 * 3.6496916e-32 = 1.9632681e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111011111011010001010111100111;
		b = 32'b10010101011011111111010011000100;
		correct = 32'b11100101111111001111000000000001;
		#400 //0.007235277 * -4.8458752e-26 = -1.4930796e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100011000001101111101000110110;
		b = 32'b00101100010000101000000111101100;
		correct = 32'b10110110001100011010011001010110;
		#400 //-7.317139e-18 * 2.764118e-12 = -2.6471876e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111111010101000111001101001110;
		b = 32'b11001011111111001000101111110010;
		correct = 32'b11110010110101110101101100000000;
		#400 //2.8239503e+38 * -33101796.0 = -8.531109e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110101110100110000001000111011;
		b = 32'b11011011111001111110100001001111;
		correct = 32'b01011001011010001110111000011100;
		#400 //-5.3497064e+32 * -1.3055229e+17 = 4097750000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100111101010111111111001111111;
		b = 32'b10110101000011100110011011001011;
		correct = 32'b01110010000110101001100110001100;
		#400 //-1.6244386e+24 * -5.3048706e-07 = 3.0621644e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101100010001101001101110101101;
		b = 32'b00001111010110011111011010001001;
		correct = 32'b11011100011010010100010001110110;
		#400 //-2.822391e-12 * 1.0746407e-29 = -2.6263577e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100110001011000100000100010011;
		b = 32'b10111010101011111110111101100010;
		correct = 32'b00101010111110101010010011011101;
		#400 //-5.976268e-16 * -0.0013422782 = 4.4523318e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010101011111110000110111010101;
		b = 32'b10111100111000111010100110000111;
		correct = 32'b00011000000011110110011010010011;
		#400 //-5.150775e-26 * -0.027790798 = 1.8534104e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110111010100101110101100000001;
		b = 32'b01101001001000001011101010111101;
		correct = 32'b00001101101001111111011111110111;
		#400 //1.25716915e-05 * 1.2144374e+25 = 1.0351865e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000110001001111001100100000111;
		b = 32'b00010001101101010000100000110111;
		correct = 32'b11110011111011010000000010011001;
		#400 //-10726.257 * 2.8561828e-28 = -3.755452e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110001010100100001101011110101;
		b = 32'b00110011101000111001110101000101;
		correct = 32'b01111101001001000101111100000101;
		#400 //1.04039106e+30 * 7.618886e-08 = 1.3655423e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011001100010010000000100001111;
		b = 32'b10100101011001100110001010111010;
		correct = 32'b00110011100110000011110001111110;
		#400 //-1.4165896e-23 * -1.998277e-16 = 7.089055e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111101100101100110110010010000;
		b = 32'b00000100100100011101101110101100;
		correct = 32'b01111000100001000000000111000111;
		#400 //0.073449254 * 3.4291073e-36 = 2.141935e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000100001000011001000101101101;
		b = 32'b00010101011011000101100110111111;
		correct = 32'b00101110001011110000000000010101;
		#400 //1.8992235e-36 * 4.7730618e-26 = 3.9790466e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010110111001101110010110011011;
		b = 32'b11100000101001101111001111000000;
		correct = 32'b00110101101100010000011010001101;
		#400 //-126936910000000.0 * -9.624136e+19 = 1.3189434e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000010100100101100101101111110;
		b = 32'b10001010110110010010101110111110;
		correct = 32'b10110111001011010000101010000111;
		#400 //2.156957e-37 * -2.0912794e-32 = -1.0314055e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001011100101111011010101001111;
		b = 32'b10011111001101011100100111100101;
		correct = 32'b00101011110101011010001111010000;
		#400 //-5.843589e-32 * -3.8495244e-20 = 1.5180027e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011100010000101010101010101001;
		b = 32'b01011010111110001010110011100011;
		correct = 32'b00000000110010000110011010000111;
		#400 //6.440979e-22 * 3.4997943e+16 = 1.8403879e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011011110001000010010101000110;
		b = 32'b00100111001001001100001100110111;
		correct = 32'b01110100000110000110000101110111;
		#400 //1.1042016e+17 * 2.2865398e-15 = 4.829138e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101001011111000000010110110011;
		b = 32'b11010000001001000011111010101101;
		correct = 32'b00011000110001000110100000110111;
		#400 //-5.5960184e-14 * -11022284000.0 = 5.0770043e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110000010101111001101010100110;
		b = 32'b10110111010011010110000010101111;
		correct = 32'b10111000100001100101111110100000;
		#400 //7.8436313e-10 * -1.2241463e-05 = -6.4074295e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001110111100101101000001101110;
		b = 32'b11101101111100001011111110011001;
		correct = 32'b00100000100000010001100100101011;
		#400 //-2036873000.0 * -9.313504e+27 = 2.1870105e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110101100100011111010110000100;
		b = 32'b01001011111100010011010110001101;
		correct = 32'b00101001000110101110100011000000;
		#400 //1.0874796e-06 * 31615770.0 = 3.4396748e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101111001110010110001000110000;
		b = 32'b11010111010100111011111010100100;
		correct = 32'b10010111011000000010000100011001;
		#400 //1.6860535e-10 * -232815750000000.0 = -7.242008e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010111101101001001011011001000;
		b = 32'b01100111000001110010001001010010;
		correct = 32'b00110000001010110000111000100101;
		#400 //397119400000000.0 * 6.381526e+23 = 6.222954e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111001001101110101010110000110;
		b = 32'b10001010001001101110101100100000;
		correct = 32'b11101110100011001001011010010011;
		#400 //0.000174841 * -8.036831e-33 = -2.1754967e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100111011001011100011010000010;
		b = 32'b01000010100010000010111101110001;
		correct = 32'b00100100010101111111011100000110;
		#400 //3.1887745e-15 * 68.09266 = 4.682993e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110101011110000101010011111111;
		b = 32'b01010111111100100101111100001110;
		correct = 32'b00011101000000110010010111011111;
		#400 //9.2510885e-07 * 532980140000000.0 = 1.7357285e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001111110100111101011001010011;
		b = 32'b10111110100100011010011111110011;
		correct = 32'b10010000101110100010100010101010;
		#400 //2.0888761e-29 * -0.28448448 = -7.342672e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111001111001011001111100001001;
		b = 32'b11001001011100111010010000001101;
		correct = 32'b11101111111100010100010011101101;
		#400 //1.490327e+35 * -997952.8 = -1.4933843e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100000100010110111000101000110;
		b = 32'b01100111111100100100101100100001;
		correct = 32'b00111000000100110101010010101011;
		#400 //8.038311e+19 * 2.2883971e+24 = 3.5126384e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101111010101110110000000100101;
		b = 32'b01000001110110000010111001110110;
		correct = 32'b11101100111111110000101110101111;
		#400 //-6.665551e+28 * 27.022686 = -2.46665e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100000011000001101001011110101;
		b = 32'b01101000100101111110100111011011;
		correct = 32'b00110111001111010110111011101110;
		#400 //6.480112e+19 * 5.7391297e+24 = 1.1291106e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100110000000101010001000000000;
		b = 32'b01110101101010111111010000001010;
		correct = 32'b10101111110000100111101110101010;
		#400 //-1.54224e+23 * 4.3595335e+32 = -3.5376263e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101001100100110111010000011000;
		b = 32'b01110001011111101010111001000000;
		correct = 32'b10110111100101000011011110100100;
		#400 //-2.2282542e+25 * 1.2611176e+30 = -1.7668885e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111111000100101111110111000100;
		b = 32'b11010100011101100111000010011101;
		correct = 32'b10101010000110001011000110001000;
		#400 //0.57418466 * -4233805200000.0 = -1.3561906e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101011010100010111110111010110;
		b = 32'b01001010001000010011011000110000;
		correct = 32'b00100000101001100101010101100111;
		#400 //7.442635e-13 * 2641292.0 = 2.8178008e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101011111011010001001110101000;
		b = 32'b11111010111101010010110001110011;
		correct = 32'b10110000011101111000101110101101;
		#400 //5.732165e+26 * -6.3650713e+35 = -9.005657e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001111011010001001000110111111;
		b = 32'b11110011010011000001110011001110;
		correct = 32'b00011011100100011101100001101101;
		#400 //-3901865700.0 * -1.617146e+31 = 2.41281e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101000100011000001001101011000;
		b = 32'b00101010100010010101110101110000;
		correct = 32'b00111101100000101000011010011001;
		#400 //1.5551511e-14 * 2.4400924e-13 = 0.06373329
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101010011101101000101100000110;
		b = 32'b10100100010001111111001101101001;
		correct = 32'b11000101100111011101001110001101;
		#400 //2.1897423e-13 * -4.3357423e-17 = -5050.444
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001110011100001000010001100001;
		b = 32'b00100011100110100010110110001010;
		correct = 32'b01101010010001111010110111111111;
		#400 //1008801860.0 * 1.6716e-17 = 6.034948e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001101100110110011100101101101;
		b = 32'b00010000000011000000010011111000;
		correct = 32'b10111101000011011110011001010011;
		#400 //-9.566437e-31 * 2.761396e-29 = -0.034643482
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100110111111100101011010011110;
		b = 32'b11000101001111110000001001101001;
		correct = 32'b11100001001010100111000000110001;
		#400 //6.0053945e+23 * -3056.1506 = -1.9650192e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001111001111010011011001010001;
		b = 32'b11000001001011111111110100100100;
		correct = 32'b00001101100010011001111000011010;
		#400 //-9.3288804e-30 * -10.999302 = 8.481338e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001110100011000000010110000111;
		b = 32'b01000011100100111110110001000100;
		correct = 32'b11001010011100100101001101100011;
		#400 //-1174586200.0 * 295.84583 = -3970264.8
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111010100000101100010111011111;
		b = 32'b01000110101000000101011101100101;
		correct = 32'b01110011010100001100101010001100;
		#400 //3.3950595e+35 * 20523.697 = 1.6542143e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010000111110100110011011110000;
		b = 32'b01110001111110011011100100001101;
		correct = 32'b10011110100000000101100100100001;
		#400 //-33608400000.0 * 2.4731354e+30 = -1.358939e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011100110001111101110011010011;
		b = 32'b10100111101000010101101010111001;
		correct = 32'b01110100100111101000110001001001;
		#400 //-4.5005055e+17 * -4.478484e-15 = 1.0049173e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010111000100111100000000011110;
		b = 32'b01000001011101010010011110100000;
		correct = 32'b11010101000110100100100101100100;
		#400 //-162453350000000.0 * 15.322174 = -10602500000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010010010001010100111001001011;
		b = 32'b01011010101000011000010010110011;
		correct = 32'b10110111000111000101110001100000;
		#400 //-211855520000.0 * 2.2731688e+16 = -9.319832e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101111011000110010010010011111;
		b = 32'b00010100001111111011110000100011;
		correct = 32'b01011010100101111010001101011000;
		#400 //2.065854e-10 * 9.680139e-27 = 2.134116e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100111100110011110101110111010;
		b = 32'b10110110011011111110000110101100;
		correct = 32'b10110000101001000100001101100110;
		#400 //4.2721606e-15 * -3.5745134e-06 = -1.1951726e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000011010100001011110011001001;
		b = 32'b00111100010100100010110001010111;
		correct = 32'b00000110011111100100000001001101;
		#400 //6.134242e-37 * 0.012827954 = 4.781933e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111001110010110110100111100;
		b = 32'b00101100010101010010111110101001;
		correct = 32'b11001010010111101010101001100111;
		#400 //-1.1052292e-05 * 3.0295577e-12 = -3648153.8
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100100000100011101110010000000;
		b = 32'b00101010100000101111011010110101;
		correct = 32'b11111001000011101000111101111101;
		#400 //-1.0762666e+22 * 2.3263826e-13 = -4.626353e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110000100111010001011111100101;
		b = 32'b01000011100011000011010001011000;
		correct = 32'b00101100100011110110101100110010;
		#400 //1.1430045e-09 * 280.40894 = 4.0762055e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100111110010100101011011000000;
		b = 32'b00110010001100111100011101101001;
		correct = 32'b01110101000100000000111111110101;
		#400 //1.9110366e+24 * 1.0464512e-08 = 1.826207e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100101011111000110110001111110;
		b = 32'b00110100100010011101001001101111;
		correct = 32'b00110000011010100110111101000010;
		#400 //2.1894274e-16 * 2.567135e-07 = 8.528681e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011101100000100110000101100001;
		b = 32'b10110001110011100001101101011110;
		correct = 32'b01101011001000011111000100101100;
		#400 //-1.1743621e+18 * -5.9985004e-09 = 1.9577596e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100001100001101100111000001101;
		b = 32'b01110110011001011111101100100111;
		correct = 32'b10101010100101100000111001011010;
		#400 //-3.108389e+20 * 1.1661425e+33 = -2.665531e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111101101100000111010000001010;
		b = 32'b00001100000101111010011010001001;
		correct = 32'b01110001000101001110111101000110;
		#400 //0.08615883 * 1.1682732e-31 = 7.374887e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110011100110111110011011110101;
		b = 32'b11101111101100111111000000011111;
		correct = 32'b01000011010111011100110111010001;
		#400 //-2.4703686e+31 * -1.1137621e+29 = 221.80397
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110110100111111000110111001101;
		b = 32'b01110010111110011110100101000010;
		correct = 32'b00000011001000110111000011111000;
		#400 //4.755077e-06 * 9.900001e+30 = 4.8031077e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101100110000100011010110010111;
		b = 32'b10000111000100100010110011100110;
		correct = 32'b01100101001010100000111110111010;
		#400 //-5.5197613e-12 * -1.0997014e-34 = 5.0193275e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100111111001010000001111110001;
		b = 32'b00101010010110101100001101011010;
		correct = 32'b00111101000001011111111110101011;
		#400 //6.356454e-15 * 1.9430066e-13 = 0.032714527
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110111011001010110100100101000;
		b = 32'b11010011000011010101100011000100;
		correct = 32'b01100011110011111011111110100000;
		#400 //-4.653003e+33 * -607079600000.0 = 7.664568e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111100111100111101000001100001;
		b = 32'b00001101001001010110011100100100;
		correct = 32'b11101111001111001010111000001001;
		#400 //-0.029762449 * 5.09687e-31 = -5.8393577e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001101011111010001101001001010;
		b = 32'b01100000111111011110010011000101;
		correct = 32'b10101011111111110011001111010111;
		#400 //-265397400.0 * 1.4635971e+20 = -1.8133228e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010000111101000001101010010001;
		b = 32'b00010110000101110111000010001000;
		correct = 32'b01111010010011100101001001100000;
		#400 //32763054000.0 * 1.2233191e-25 = 2.6782098e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100100110100100111111000000011;
		b = 32'b01111011010001010000001000011101;
		correct = 32'b00101001000010001100001011000100;
		#400 //3.106317e+22 * 1.02292534e+36 = 3.0367e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011111110001011111100000010100;
		b = 32'b10101001100110011000100000001000;
		correct = 32'b00110101101001010000110001000111;
		#400 //-8.3843156e-20 * -6.8181626e-14 = 1.2297031e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111111010010001110001111110110;
		b = 32'b11000110011100000010001011000000;
		correct = 32'b01111000010101100010100101111100;
		#400 //-2.6702924e+38 * -15368.6875 = 1.737489e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000110000100111001101001000110;
		b = 32'b11000100101111111001001101101110;
		correct = 32'b00000000110001010011110100111011;
		#400 //-2.776097e-35 * -1532.6072 = 1.8113558e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010111011001101110001110011110;
		b = 32'b00000111101000100010101000111000;
		correct = 32'b11001111001101100011111011010010;
		#400 //-7.46043e-25 * 2.4399865e-34 = -3057570300.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001100110101000100110101111011;
		b = 32'b10101010100111110000000101111100;
		correct = 32'b10100001101010101110011101110010;
		#400 //3.2710404e-31 * -2.8245104e-13 = -1.1580911e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110001001011010000111101110111;
		b = 32'b11110001000011011000001000100101;
		correct = 32'b10111111100111001000101001000011;
		#400 //8.5695364e+29 * -7.0071554e+29 = -1.2229694
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000001110010011001011000010010;
		b = 32'b11010010110011010111000010011111;
		correct = 32'b10101110011110110011001010100111;
		#400 //25.198277 * -441178880000.0 = -5.711578e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101101000011010011111001010010;
		b = 32'b00111111000101010010111001011110;
		correct = 32'b01101101011100100110000011110000;
		#400 //2.7320454e+27 * 0.58273876 = 4.6882852e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111100111110101000101111010111;
		b = 32'b10000110110111101101100011011010;
		correct = 32'b01110101100011111110100011110101;
		#400 //-0.030584259 * -8.3825753e-35 = 3.6485517e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001110001010100011001110111111;
		b = 32'b00100011101011010101000011001100;
		correct = 32'b11101001111110110110011010110010;
		#400 //-713879500.0 * 1.8790916e-17 = -3.7990668e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110010110000100011010011001001;
		b = 32'b11011001100110001000011011101100;
		correct = 32'b00011000101000101111101000011010;
		#400 //-2.2608576e-08 * -5366568000000000.0 = 4.2128557e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111000100011010100000010101111;
		b = 32'b10001111000001010000110000010011;
		correct = 32'b11101001000001111110010011101100;
		#400 //6.735452e-05 * -6.559732e-30 = -1.0267877e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001101000000000001000101010101;
		b = 32'b10010011001001101000100011011101;
		correct = 32'b11111001010001001101111000110011;
		#400 //134288720.0 * -2.1019624e-27 = -6.3887307e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011000100010011000111100111010;
		b = 32'b10100001101001100100000001011010;
		correct = 32'b00110110010100111101000110110101;
		#400 //-3.555829e-24 * -1.1265631e-18 = 3.1563516e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100011101100101101001010110011;
		b = 32'b11010100001011011011101000110111;
		correct = 32'b10001111000000111100000100100000;
		#400 //1.9388033e-17 * -2984614000000.0 = -6.495993e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100011010011101101111010111000;
		b = 32'b11110001000111100000010110010001;
		correct = 32'b00110001101001111001000101011101;
		#400 //-3.8160779e+21 * -7.824858e+29 = 4.8768656e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110110110010101101100100010000;
		b = 32'b01100010101111011100000101111011;
		correct = 32'b11010011100010001101010011010000;
		#400 //-2.0571221e+33 * 1.7501882e+21 = -1175371900000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101111000101011000000100110000;
		b = 32'b01010110011100001110000001110010;
		correct = 32'b01011000000111101110010000100100;
		#400 //4.6269445e+28 * 66211694000000.0 = 698810800000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000110100001110010101110110101;
		b = 32'b00100010111001000110100100001001;
		correct = 32'b11100011000101110111111101111110;
		#400 //-17301.854 * 6.1910734e-18 = -2.794645e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111100101001100110101011110110;
		b = 32'b11001000000101100110000100001110;
		correct = 32'b11110100000011011010011011100000;
		#400 //6.9127256e+36 * -153988.22 = -4.4891265e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011010011101110000110110011010;
		b = 32'b11001001001000000010011001010001;
		correct = 32'b11010000110001010111010100110010;
		#400 //1.7384819e+16 * -655973.06 = -26502337000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101001101001010100111001000111;
		b = 32'b11010110111110110010010000001011;
		correct = 32'b11010010001010001000000100010011;
		#400 //2.4980302e+25 * -138066110000000.0 = -180930000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100110000001100110011101010011;
		b = 32'b11111111000010111111111101110010;
		correct = 32'b10100110011101011100010100111001;
		#400 //1.5867578e+23 * -1.8608904e+38 = -8.5268737e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101000100001000010100010010000;
		b = 32'b01011100011011111110011011111111;
		correct = 32'b11001011100011010000011011000010;
		#400 //-4.992805e+24 * 2.7010601e+17 = -18484612.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010111111111010110001111101110;
		b = 32'b01010110000010101111100101111000;
		correct = 32'b11000001011010010110000101110110;
		#400 //-557211270000000.0 * 38201016000000.0 = -14.586294
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010111111101101101100111101010;
		b = 32'b10110101010101110100000001000010;
		correct = 32'b11100010000100101100101010001101;
		#400 //542831600000000.0 * -8.018725e-07 = -6.76955e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101110100010000101100101111100;
		b = 32'b01011001011100000111110110011111;
		correct = 32'b10010100100100010010010010001100;
		#400 //-6.2004596e-11 * 4230757300000000.0 = -1.4655674e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011000000001100010111110011000;
		b = 32'b01011000011011010000011111001110;
		correct = 32'b00111111000100001110110010111111;
		#400 //590155900000000.0 * 1042471100000000.0 = 0.56611246
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100011101011010110100001111010;
		b = 32'b01111101000111111101011010011010;
		correct = 32'b10100110000010101101110111101001;
		#400 //-6.39763e+21 * 1.3278845e+37 = -4.817911e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110101101011111110000110010;
		b = 32'b01101101011111000010101100100001;
		correct = 32'b00010000101110001100000000010010;
		#400 //0.35543972 * 4.8776476e+27 = 7.2871134e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110011001100001001001010111000;
		b = 32'b10110111010000110010101001000100;
		correct = 32'b00111011011001111001110011011011;
		#400 //-4.1111633e-08 * -1.16327465e-05 = 0.0035341296
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101000101000000001101110000001;
		b = 32'b10010000111000110111000010000100;
		correct = 32'b11010111001101000011011001111000;
		#400 //1.7775496e-14 * -8.970907e-29 = -198146030000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001111001101110010111100101000;
		b = 32'b01010000000100111001001101101101;
		correct = 32'b10111110100111101110001010001000;
		#400 //-3073321000.0 * 9903650000.0 = -0.31032205
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011110101000101110000111100100;
		b = 32'b00111101000001101101011011001000;
		correct = 32'b11100001000110101001111011111101;
		#400 //-5.8684564e+18 * 0.032919675 = -1.7826593e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111100110100110100010001011010;
		b = 32'b01001101000001000001110110110010;
		correct = 32'b01101111010011001010111101100011;
		#400 //8.775688e+36 * 138533660.0 = 6.334697e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100111011010101001010101100001;
		b = 32'b10110111110101100100011000000110;
		correct = 32'b01101111000011000010000111101101;
		#400 //-1.1077893e+24 * -2.5543395e-05 = 4.3368915e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100010000011010000110000100111;
		b = 32'b00100010101110110001100000101111;
		correct = 32'b01111110110000001111111010000110;
		#400 //6.5046665e+20 * 5.0712057e-18 = 1.2826667e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010000000111110010011101001010;
		b = 32'b00111101010001011111101011100000;
		correct = 32'b00010010010011011100101110000101;
		#400 //3.1387488e-29 * 0.048334956 = 6.493745e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011111100110100011011001001111;
		b = 32'b10101001111110010011011000000000;
		correct = 32'b11110101000111100110100111001001;
		#400 //2.2224312e+19 * -1.1067189e-13 = -2.0081262e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010110000000111010100100011100;
		b = 32'b00110011000000010000100011111000;
		correct = 32'b01100010100000101001101011000000;
		#400 //36190586000000.0 * 3.004331e-08 = 1.2046138e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110000000110111010010111011100;
		b = 32'b11000100010011001100011001001100;
		correct = 32'b01101011010000101001010110000001;
		#400 //-1.9268275e+29 * -819.0984 = 2.3523762e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010000111001001000110010001010;
		b = 32'b11000001110111100101100110100011;
		correct = 32'b11001110100000111001000110001000;
		#400 //30675325000.0 * -27.793768 = -1103676400.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010000110010011011101010110100;
		b = 32'b00111000101011001001100101110010;
		correct = 32'b00010111100101011001101001010001;
		#400 //7.956818e-29 * 8.2301805e-05 = 9.667854e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101001101101011010010101100111;
		b = 32'b11001001001100101000011101011010;
		correct = 32'b00100000000000100011110000101110;
		#400 //-8.0667074e-14 * -731253.6 = 1.103134e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000010101110010010011000011000;
		b = 32'b11110111010110010011011000101101;
		correct = 32'b00001010110110100011011000101011;
		#400 //-92.5744 * -4.405575e+33 = 2.1013012e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000101001001100101111011101100;
		b = 32'b10101001111101100100111101001000;
		correct = 32'b01011010101011001110101010001000;
		#400 //-2661.9326 * -1.0938348e-13 = 2.4335783e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010011100000011110001110101000;
		b = 32'b11001001010001001000000001010011;
		correct = 32'b01001001101010010011011111110010;
		#400 //-1115740400000.0 * -804869.2 = 1386238.2
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101110001111101011100101100110;
		b = 32'b01100110000000101100000110001010;
		correct = 32'b00000111101110101011010001001000;
		#400 //4.3365665e-11 * 1.5436945e+23 = 2.809213e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111000111111000101011100101;
		b = 32'b00010110101000001010001110011010;
		correct = 32'b11011111111111100100000010101000;
		#400 //-9.509477e-06 * 2.5952641e-25 = -3.6641656e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011111011011100101011100001111;
		b = 32'b10101110000011000011110000010010;
		correct = 32'b00110000110110011000101111011010;
		#400 //-5.0470474e-20 * -3.1885668e-11 = 1.5828576e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100110010100010101111001011110;
		b = 32'b01101001110001100111101110000000;
		correct = 32'b00111100000001110000010100111011;
		#400 //2.4717884e+23 * 2.9993816e+25 = 0.008240993
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101011001010011010001000100011;
		b = 32'b11011111000010100001000000010100;
		correct = 32'b10001011100111010100010011111110;
		#400 //6.026587e-13 * -9.948474e+18 = -6.057801e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101001000000101010001011001100;
		b = 32'b00100011001110101011011100000110;
		correct = 32'b11000101001100110001110010001101;
		#400 //-2.9007002e-14 * 1.0121837e-17 = -2865.7844
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000101010101110110000110001110;
		b = 32'b01011000101111111110111010100011;
		correct = 32'b00101100000011111010001101011100;
		#400 //3446.0972 * 1688253300000000.0 = 2.0412205e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011101100111100100010101111111;
		b = 32'b10101111101101011001010111101001;
		correct = 32'b11101101010111110010000110110101;
		#400 //1.4255827e+18 * -3.3030226e-10 = -4.3159942e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100111011000010100011010110110;
		b = 32'b11000101001001110110110010101000;
		correct = 32'b10100001101011000011101010100100;
		#400 //3.1263355e-15 * -2678.791 = -1.1670695e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110011000110101011111011100100;
		b = 32'b01010110000100101111100011110111;
		correct = 32'b00011100100001101100010100001100;
		#400 //3.6029533e-08 * 40399500000000.0 = 8.918312e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110101111110110101000010110101;
		b = 32'b11011111101111011001110011011000;
		correct = 32'b10010101101010011010011100101001;
		#400 //1.8724446e-06 * -2.7326066e+19 = -6.852229e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110010011000011011000111111000;
		b = 32'b10111001100100111111111010010111;
		correct = 32'b00111000010000110011001111111111;
		#400 //-1.3137189e-08 * -0.0002822771 = 4.6540048e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110110011110001110111101111000;
		b = 32'b01101110101010000110111000011001;
		correct = 32'b01000111001111010010111001001001;
		#400 //1.2622526e+33 * 2.606329e+28 = 48430.285
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110100010011110010111100000001;
		b = 32'b11000001010110101011110111001010;
		correct = 32'b10110010011100100111100100111101;
		#400 //1.9295477e-07 * -13.671335 = -1.411382e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000001111111001000001110001100;
		b = 32'b10110011111001011110110010011111;
		correct = 32'b01001101100011001001001101100010;
		#400 //-31.564232 * -1.07066846e-07 = 294808640.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001111001100010000010101010111;
		b = 32'b00110010111100010101000000100101;
		correct = 32'b10011011101110111100101101111000;
		#400 //-8.727802e-30 * 2.8092538e-08 = -3.1068044e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110101110000100010000010110100;
		b = 32'b01001101010111000001110101001001;
		correct = 32'b10100111111000011100011011010110;
		#400 //-1.4463644e-06 * 230806670.0 = -6.2665623e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100010100011011110010111111001;
		b = 32'b11011010100110101001011100100011;
		correct = 32'b01000111011010101111101101101011;
		#400 //-1.3087811e+21 * -2.1756661e+16 = 60155.418
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001010011110001011101011110001;
		b = 32'b11101101011100001101010000101011;
		correct = 32'b10011100100001000011001100011010;
		#400 //4075196.2 * -4.658306e+27 = -8.748237e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010010011010011100000010000111;
		b = 32'b10111111101001111000101000010101;
		correct = 32'b10010010001100101001011000100010;
		#400 //7.3759145e-28 * -1.3089014 = -5.635195e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011001001110100000010100011111;
		b = 32'b11001000001100110000000100010111;
		correct = 32'b00010000100001010000010001001000;
		#400 //-9.617009e-24 * -183300.36 = 5.2465847e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011010110101100110110011000101;
		b = 32'b00100001101100111110010010101101;
		correct = 32'b10111000100110001001001000000101;
		#400 //-8.868405e-23 * 1.2190042e-18 = -7.275123e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000100000100000100111110100000;
		b = 32'b00100000000011001101001010111110;
		correct = 32'b11100011100000110010101110010100;
		#400 //-577.24414 * 1.192819e-19 = -4.839327e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010110011111111101001110001001;
		b = 32'b10001111010010000100110011000001;
		correct = 32'b11000110101000110111101111011000;
		#400 //2.0665485e-25 * -9.8755436e-30 = -20925.922
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110001101011111001101000101000;
		b = 32'b00110111011101101001110000111010;
		correct = 32'b01111001101101100100100111001100;
		#400 //1.7390797e+30 * 1.4699117e-05 = 1.1831185e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000011101011010110110101010011;
		b = 32'b11110111111101000110011111001010;
		correct = 32'b00001011001101011010011110001000;
		#400 //-346.8541 * -9.914262e+33 = 3.4985368e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010110100111011110000101100010;
		b = 32'b00000101111101000101010001111000;
		correct = 32'b01010000001001010110101111011011;
		#400 //2.5506955e-25 * 2.2976679e-35 = 11101236000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000101001101011000100100001110;
		b = 32'b00011110000000111010111001011101;
		correct = 32'b10100110101100000111010111101010;
		#400 //-8.535752e-36 * 6.97114e-21 = -1.2244414e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010010000101100101101011010010;
		b = 32'b00110100101010011110111001111000;
		correct = 32'b11011100111000101000001000000001;
		#400 //-161442200000.0 * 3.1652212e-07 = -5.100503e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000010100010000001110101000110;
		b = 32'b00101111011111101100100010100111;
		correct = 32'b10010010100010001100001110011011;
		#400 //-2.0000206e-37 * 2.3172451e-10 = -8.631027e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000010110101111101110011110110;
		b = 32'b10110110010100001000100110110010;
		correct = 32'b10001100000001000111111100001000;
		#400 //3.1718236e-37 * -3.1074565e-06 = -1.0207137e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000100101110001000010101111;
		b = 32'b11011110010111110001111111001010;
		correct = 32'b00010001101011010101001011010111;
		#400 //-1.0991438e-09 * -4.0194478e+18 = 2.7345641e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110100001101000101011011110101;
		b = 32'b00000110101111000000111001000111;
		correct = 32'b11101100111101010111111100000000;
		#400 //-1.6795441e-07 * 7.073872e-35 = -2.3742925e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001110101111000011101010110110;
		b = 32'b10110010101000101110001111001110;
		correct = 32'b11011011100100111110100101110101;
		#400 //1578982100.0 * -1.8962876e-08 = -8.326702e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101110001001011110111011001001;
		b = 32'b01000010101011101000100100110101;
		correct = 32'b00101010111100110110000110011011;
		#400 //3.772874e-11 * 87.26798 = 4.3233199e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111111011011011111000101111110;
		b = 32'b11010000101111100001010001100010;
		correct = 32'b00101110001000000011101101000101;
		#400 //-0.9294661 * -25512055000.0 = 3.643243e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000011111000101111110110010101;
		b = 32'b10000111010000011000100010011110;
		correct = 32'b10111100000101100010000010111010;
		#400 //1.3341306e-36 * -1.4559854e-34 = -0.009163076
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111101011111110101110011000100;
		b = 32'b11110011100000010100100100110001;
		correct = 32'b00001001011111001101001010001110;
		#400 //-0.062344328 * -2.048617e+31 = 3.0432399e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111100010111100110000110110010;
		b = 32'b10010000110111001111100100100001;
		correct = 32'b01101011000000001101000011011100;
		#400 //-0.013573097 * -8.7158543e-29 = 1.5572882e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111010100001001000010011101110;
		b = 32'b11110000001110111001011010001010;
		correct = 32'b11001001101101001101100100011001;
		#400 //3.4403966e+35 * -2.3222275e+29 = -1481507.1
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011010011101000011011011001111;
		b = 32'b11000101010010101010110000100110;
		correct = 32'b10010100100110100011110001110000;
		#400 //5.050229e-23 * -3242.7593 = -1.5573865e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110111110101011101001111001010;
		b = 32'b01001110011101001000101111001111;
		correct = 32'b11101000110111111101011110100111;
		#400 //-8.673866e+33 * 1025700800.0 = -8.4565265e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101110110010111011011001100000;
		b = 32'b00101100011011111111001100001001;
		correct = 32'b01000001110110010101011011001111;
		#400 //9.2637675e-11 * 3.4098854e-12 = 27.167387
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110010101101100110101001000100;
		b = 32'b11100010010010100011011001000100;
		correct = 32'b10001111111001101110111111101100;
		#400 //2.1235913e-08 * -9.3253814e+20 = -2.2772166e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111011101100011101011101110110;
		b = 32'b00101000000100111010000101011110;
		correct = 32'b11010011000110100011000110110010;
		#400 //-0.0054272963 * 8.19513e-15 = -662258700000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101100000110110101100010111111;
		b = 32'b00111111101111100110101000001010;
		correct = 32'b10101011110100001101101010010111;
		#400 //-2.2076089e-12 * 1.487611 = -1.483996e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110111011001000110011011010101;
		b = 32'b11100101010001101001101111011111;
		correct = 32'b11010001100100110011001101110010;
		#400 //4.6325366e+33 * -5.8618992e+22 = -79027910000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001100100100110001100001001011;
		b = 32'b10010010100000101110011101101010;
		correct = 32'b01111001100011111101010011101110;
		#400 //-77120090.0 * -8.261201e-28 = 9.335215e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001000101101110000101001100010;
		b = 32'b00100101101110011010000000110010;
		correct = 32'b00100010011111000110111101001000;
		#400 //1.1016353e-33 * 3.2200937e-16 = 3.421128e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111001110011011110100000101011;
		b = 32'b11011100100100010110001110100110;
		correct = 32'b01011100101101010100011110001010;
		#400 //-1.3364122e+35 * -3.273875e+17 = 4.0820503e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110100010111010111101100101111;
		b = 32'b01110001010111110100011101000000;
		correct = 32'b11000010011111011111000010000011;
		#400 //-7.019019e+31 * 1.1056207e+30 = -63.484875
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111000110010110110010110001100;
		b = 32'b01010000110001101111000001000110;
		correct = 32'b10100111100000101101111001010000;
		#400 //-9.698709e-05 * 26701083000.0 = -3.632328e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011110110001110010110110010;
		b = 32'b11001101001110001100010001110011;
		correct = 32'b00111110000101100100001000100101;
		#400 //-28429156.0 * -193742640.0 = 0.1467367
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101100010111111000111101100000;
		b = 32'b10101101111001110001000101101100;
		correct = 32'b00111101111101111010111010010001;
		#400 //-3.1769795e-12 * -2.6269396e-11 = 0.12093843
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010011000110111100001101100000;
		b = 32'b00011010010111100011001111011011;
		correct = 32'b01111000001100110111010001111111;
		#400 //668997800000.0 * 4.5950413e-23 = 1.4559124e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111001011100011110001111111001;
		b = 32'b01001011111010011111000011010010;
		correct = 32'b11101101000001000101100110000111;
		#400 //-7.849796e+34 * 30663076.0 = -2.5600158e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111011110010011000011011111110;
		b = 32'b10101011000100000010001001000101;
		correct = 32'b01010000001100101111100000010001;
		#400 //-0.0061501255 * -5.1206636e-13 = 12010407000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011001100110110100010111001111;
		b = 32'b00000010111111111000111000100011;
		correct = 32'b01010110000110111000101011111110;
		#400 //1.605482e-23 * 3.7550465e-37 = 42755317000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110000011001111000011001111101;
		b = 32'b01011100011011101101100011001100;
		correct = 32'b00010011011110000010011100010110;
		#400 //8.422843e-10 * 2.6891766e+17 = 3.1321272e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001011011011101011100100011011;
		b = 32'b11101011001100011100011011111101;
		correct = 32'b10011111101010111110000110001110;
		#400 //15644955.0 * -2.1491957e+26 = -7.2794466e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101000110110000110011101010011;
		b = 32'b01000111011011101110000001100100;
		correct = 32'b11100000111001111110101010001001;
		#400 //-8.175497e+24 * 61152.39 = -1.3369056e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111111111110111011010000100001;
		b = 32'b01000011110001100110010011101000;
		correct = 32'b10111011101000100110010011101011;
		#400 //-1.9664346 * 396.78833 = -0.004955878
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001100110100001001101111110011;
		b = 32'b10111001010100101011111011000111;
		correct = 32'b11010010111111010110011110111111;
		#400 //109371290.0 * -0.00020098231 = -544183650000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000011111000101101011010111111;
		b = 32'b01110101011100001010111111000000;
		correct = 32'b00001101111100010100010101110011;
		#400 //453.6777 * 3.0510642e+32 = 1.4869491e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000011111000101010100001110100;
		b = 32'b10011011011011001101110010010100;
		correct = 32'b10100111111101001111100011010001;
		#400 //1.3321761e-36 * -1.9592735e-22 = -6.799337e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100010010010011110101000100011;
		b = 32'b10011101010111001101010111010010;
		correct = 32'b11000100011010100001000100001000;
		#400 //2.736453e-18 * -2.92273e-21 = -936.2661
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000011101011000110001101101110;
		b = 32'b11000010101000000000111010010100;
		correct = 32'b10000000100010011101110010010101;
		#400 //1.0132079e-36 * -80.02847 = -1.2660593e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100000001011100000100011111;
		b = 32'b00000111011100001000010001111111;
		correct = 32'b01111100000011100101110101000101;
		#400 //535.0175 * 1.809453e-34 = 2.9567915e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011011011101010001111100100111;
		b = 32'b10011110101010001011011101101000;
		correct = 32'b00111100001110011111011101100010;
		#400 //-2.0275991e-22 * -1.7863547e-20 = 0.011350485
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111010010111011010101111001100;
		b = 32'b01011111011011100011000010111000;
		correct = 32'b01011010011011100011111011100001;
		#400 //2.8774552e+35 * 1.716342e+19 = 1.6765045e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011101010010001111011001110100;
		b = 32'b10011000110001100011001100111111;
		correct = 32'b01000100000000011100100010111001;
		#400 //-2.6597193e-21 * -5.1233546e-24 = 519.1363
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011010001100000010100111000110;
		b = 32'b00110100101101100011101101101001;
		correct = 32'b10100100111101110111100101110011;
		#400 //-3.642969e-23 * 3.3943368e-07 = -1.0732492e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100110010110110010010001110011;
		b = 32'b01000001101100110111101101111101;
		correct = 32'b11100100000111000100100010110101;
		#400 //-2.5871766e+23 * 22.435297 = -1.1531725e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000100001010001100000000110000;
		b = 32'b10110111101110101100110010110110;
		correct = 32'b00001011111001110100001111001011;
		#400 //-1.9836553e-36 * -2.2268254e-05 = 8.9079967e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101101011110010000111001110011;
		b = 32'b00111101100011111011111010100101;
		correct = 32'b00101111010111011100011011010101;
		#400 //1.415722e-11 * 0.070187844 = 2.0170472e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110011000110100011001011011101;
		b = 32'b01110111100111111101111110001011;
		correct = 32'b10111010111101101110100111011111;
		#400 //-1.2216878e+31 * 6.485228e+33 = -0.001883801
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100000010100000110111100011100;
		b = 32'b10101110101010111101100111111100;
		correct = 32'b01110001000110110011111101101011;
		#400 //-6.0077016e+19 * -7.8149015e-11 = 7.687495e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010010000010011111000101111010;
		b = 32'b10100111011101010001011010001111;
		correct = 32'b01101010000100000001010110110110;
		#400 //-148115460000.0 * -3.401281e-15 = 4.354696e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001111011001000100000100011011;
		b = 32'b01010011010011010001010001001000;
		correct = 32'b00111011100011100111011011110111;
		#400 //3829472000.0 * 880808560000.0 = 0.004347678
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011010011011101001101110111100;
		b = 32'b10010001010101011101111000101010;
		correct = 32'b11001000100011101100111010100101;
		#400 //4.9343048e-23 * -1.6871197e-28 = -292469.16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010011001011010001001001010011;
		b = 32'b00001101101010111000100110100100;
		correct = 32'b11000101000000010010010100000100;
		#400 //-2.1844704e-27 * 1.0571824e-30 = -2066.3135
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111101001010010101011100110111;
		b = 32'b10000001100100011110010100111000;
		correct = 32'b01111011000101001001000111001100;
		#400 //-0.04134294 * -5.35935e-38 = 7.7141705e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000000110100000100010010000000;
		b = 32'b01010000010000101011010011101010;
		correct = 32'b00110000000010001110101000111000;
		#400 //6.508362 * 13066545000.0 = 4.9809357e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000110001000111100001100111011;
		b = 32'b01111101100010001100111010011011;
		correct = 32'b00001000000110010011100001100100;
		#400 //10480.808 * 2.273097e+37 = 4.610805e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110011111101101010111000111101;
		b = 32'b11010111000001101001011011011010;
		correct = 32'b10011100011010101001101010000010;
		#400 //1.14869614e-07 * -147982460000000.0 = -7.76238e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101110010101111100110010000110;
		b = 32'b01001001001000111011101100111111;
		correct = 32'b10100100101010001011010001100111;
		#400 //-4.9066994e-11 * 670643.94 = -7.3164e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111111011011000101011001001011;
		b = 32'b11001010001000101101101100110000;
		correct = 32'b11110100101110011100000011110100;
		#400 //3.1414587e+38 * -2668236.0 = -1.1773541e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110101010011001001011100100001;
		b = 32'b01110110000110111100011011010011;
		correct = 32'b10111110101010000001110000010100;
		#400 //-2.5934908e+32 * 7.898815e+32 = -0.32833922
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000100000000111101111111101011;
		b = 32'b01001000010010011000111101110001;
		correct = 32'b10111011001001110111111000101101;
		#400 //-527.4987 * 206397.77 = -0.0025557384
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010001101100111101101110010001;
		b = 32'b10011001101100101100111000101011;
		correct = 32'b01110111100000001100000011011010;
		#400 //-96560360000.0 * -1.8488039e-23 = 5.2228554e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100001110000010111000001110101;
		b = 32'b01111010000011101010010010111011;
		correct = 32'b10100111001011011001010011001011;
		#400 //-4.4604062e+20 * 1.8516182e+35 = -2.4089234e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100110001001110110001111010;
		b = 32'b00011101000000101110010110110111;
		correct = 32'b01100111010000001001000010100001;
		#400 //1575.3899 * 1.7324117e-21 = 9.093623e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100111110000110011111110100101;
		b = 32'b11100101100000000011000000101111;
		correct = 32'b10000001110000101111011001000001;
		#400 //5.4192376e-15 * -7.566897e+22 = -7.16177e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010100100111100001001101000010;
		b = 32'b00111011001000111111001000101010;
		correct = 32'b01011000111101101101010100111010;
		#400 //5431423400000.0 * 0.0025016167 = 2171165300000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111011100101000001100011101100;
		b = 32'b00111110100100100011110110101110;
		correct = 32'b11111100100000011001111111110111;
		#400 //-1.5379308e+36 * 0.28562683 = -5.384406e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110110010111111000001000000100;
		b = 32'b00111111011011101111001110011110;
		correct = 32'b00110110011011110111010001010011;
		#400 //3.3305269e-06 * 0.9334048 = 3.5681485e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010011001100001010000011101100;
		b = 32'b11101001110111010010011111100101;
		correct = 32'b00101000110011000111010100010001;
		#400 //-758614070000.0 * -3.3420125e+25 = 2.269932e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001000110100011001110001010110;
		b = 32'b01001001110100100010101101000101;
		correct = 32'b00111110011111110101000111100110;
		#400 //429282.7 * 1721704.6 = 0.24933586
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101000001110010011011111010000;
		b = 32'b10110111101110100010111011001100;
		correct = 32'b10101111111111101010110001100110;
		#400 //1.0281665e-14 * -2.219472e-05 = -4.6324827e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010000000110110010100000001111;
		b = 32'b11101010000100100001010011111110;
		correct = 32'b10100101100001111111001110000101;
		#400 //10412375000.0 * -4.4150576e+25 = -2.3583782e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111101010000100010110001000001;
		b = 32'b10001110001011110011101001010011;
		correct = 32'b11101110100011011101011011000100;
		#400 //0.047405485 * -2.1598497e-30 = -2.194851e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101000010100100111101010000110;
		b = 32'b00001110010111001000110110100000;
		correct = 32'b01011001011101000100111001100100;
		#400 //1.168391e-14 * 2.7185284e-30 = 4297880400000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001100000110011110101100000010;
		b = 32'b01111100011100100000111100110110;
		correct = 32'b10001111001000101100100001001010;
		#400 //-40348680.0 * 5.0273774e+36 = -8.025791e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101000101001010001110001101010;
		b = 32'b00111000011111111010110010100011;
		correct = 32'b00101111101001010101001001000000;
		#400 //1.8331003e-14 * 6.0957518e-05 = 3.0071767e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000011010010101010111010001110;
		b = 32'b00011110100101111101100001101011;
		correct = 32'b01100100001010101101101001101111;
		#400 //202.68185 * 1.6077255e-20 = 1.2606745e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110000111011011110111100111001;
		b = 32'b01000011110101001010000100111010;
		correct = 32'b00101100100011110011101110101000;
		#400 //1.7312011e-09 * 425.25958 = 4.0709276e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100110110011011111010011010010;
		b = 32'b01011000100000101010001111101111;
		correct = 32'b11001101110010011100101100110100;
		#400 //-4.8630063e+23 * 1149124800000000.0 = -423192200.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110111101101000100001011110110;
		b = 32'b11011101000011110110010001010110;
		correct = 32'b10011010001000001110100101110111;
		#400 //2.1488853e-05 * -6.457799e+17 = -3.3275816e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110001110101100000111100100001;
		b = 32'b01010100111100010101001000111101;
		correct = 32'b01011100011000110001010001100000;
		#400 //2.1199386e+30 * 8291735000000.0 = 2.5566889e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001100011000011000000100100111;
		b = 32'b00000101011110111000110101000010;
		correct = 32'b11000110011001010111110111111011;
		#400 //-1.7372235e-31 * 1.1827908e-35 = -14687.495
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001000000000010001110110011101;
		b = 32'b11010111100110010101001100010000;
		correct = 32'b00101111110101111001010001011011;
		#400 //-132214.45 * -337164060000000.0 = 3.9213685e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001010001000110111000110001100;
		b = 32'b01011101010111101010010000010000;
		correct = 32'b00101100001110111110111011010011;
		#400 //2677859.0 * 1.00268534e+18 = 2.6706872e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111001000001111011100011001101;
		b = 32'b01111000011011000011001001010000;
		correct = 32'b11000000000100110001100111101010;
		#400 //-4.404427e+34 * 1.9162539e+34 = -2.2984567
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010001000100010101001100010;
		b = 32'b01101111011111001101000110100010;
		correct = 32'b10001010001001000011010010111110;
		#400 //-0.0006186125 * 7.8243653e+28 = -7.9062325e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001011011011001000101111000001;
		b = 32'b10001110001111101101101011101011;
		correct = 32'b11111100100111101010010010101011;
		#400 //15502273.0 * -2.3524713e-30 = -6.589782e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010010110011001011011100011011;
		b = 32'b11000001001100000100011010100011;
		correct = 32'b01010001000101001010011010011001;
		#400 //-439622660000.0 * -11.017245 = 39903138000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110011111100101100101011011100;
		b = 32'b11011110111100101010100000110000;
		correct = 32'b01010100100000000001001001001010;
		#400 //-3.8471995e+31 * -8.742639e+18 = 4400501000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110111011001011110110010100001;
		b = 32'b11110011111101100100101110101000;
		correct = 32'b11000010111011101111101111010111;
		#400 //4.6634195e+33 * -3.9027085e+31 = -119.491875
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010110101010100111101110010011;
		b = 32'b01001001001011001101101101100101;
		correct = 32'b10001100111111000111101111010011;
		#400 //-2.7542968e-25 * 708022.3 = -3.8901272e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010001110100000110001001010011;
		b = 32'b00011110011000011010111010000101;
		correct = 32'b10110010111011000110000011101011;
		#400 //-3.287721e-28 * 1.1947491e-20 = -2.751809e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101001100110001010001010011111;
		b = 32'b11010010111101000010111101001000;
		correct = 32'b01010110001000000000010101010001;
		#400 //-2.3065585e+25 * -524382630000.0 = 43986174000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010011100010011111000001010010;
		b = 32'b10001111000011010001001011000011;
		correct = 32'b01000011111110100100111111011000;
		#400 //-3.4820636e-27 * -6.95545e-30 = 500.62378
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101000010110001011011010001111;
		b = 32'b10011001111001010001000111010001;
		correct = 32'b01001101111100100011000011011011;
		#400 //-1.2029995e-14 * -2.3685241e-23 = 507911000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100110000110111101101011101100;
		b = 32'b01000101101001010011101000001011;
		correct = 32'b00011111111100010111101011010110;
		#400 //5.407312e-16 * 5287.2554 = 1.02270685e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101101101101010101110011000100;
		b = 32'b01001010011101110111011011000101;
		correct = 32'b11100010101110111001111001001001;
		#400 //-7.0161167e+27 * 4054449.2 = -1.7304734e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001111110000010101010111100010;
		b = 32'b01111001111010011011001110111000;
		correct = 32'b10010101010100111100100000110001;
		#400 //-6487262000.0 * 1.5168129e+35 = -4.2769034e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011011110110011110001010110001;
		b = 32'b00111011000100000010100110001000;
		correct = 32'b01100000010000010111010101000011;
		#400 //1.2265864e+17 * 0.002199741 = 5.5760488e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000011010110000110101010100100;
		b = 32'b10000111001010000000001111010101;
		correct = 32'b00111011101001001101111111000110;
		#400 //-6.3599112e-37 * -1.2640041e-34 = 0.0050315587
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010000100101100010010001110111;
		b = 32'b01001010001100101010110011111000;
		correct = 32'b11000101110101110001111001011111;
		#400 //-20151777000.0 * 2927422.0 = -6883.7964
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011010001110010110111000110001;
		b = 32'b11001010011000001011011100010010;
		correct = 32'b10001111010100110011111100000000;
		#400 //3.8346115e-23 * -3681732.5 = -1.04152365e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100000000101000101110110001100;
		b = 32'b10011000010100101101100101000110;
		correct = 32'b01000111001101000010001011110000;
		#400 //-1.256704e-19 * -2.7251559e-24 = 46114.938
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111001000110100111001010010000;
		b = 32'b00100101010011111100001010011101;
		correct = 32'b11010011001111100100111100000011;
		#400 //-0.00014729262 * 1.8020326e-16 = -817369400000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000110010100001110001111011011;
		b = 32'b00010100000100010111100101110001;
		correct = 32'b11110001101101111100110001010110;
		#400 //-13368.964 * 7.344579e-27 = -1.8202491e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100111100101101010101000010100;
		b = 32'b01000011101000010110100000100000;
		correct = 32'b01100011011011101111011001000110;
		#400 //1.4229847e+24 * 322.81348 = 4.408071e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000101100101110110100011010010;
		b = 32'b10010110000111000100110001011011;
		correct = 32'b00101110111101111111111000011110;
		#400 //-1.4238477e-35 * -1.2625673e-25 = 1.12774e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010101111111110100110001001111;
		b = 32'b11100010000100011111100110010000;
		correct = 32'b10110011010111111101110010001101;
		#400 //35087900000000.0 * -6.731902e+20 = -5.2121823e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000111011011100001110111101001;
		b = 32'b00111001010001001100111101100001;
		correct = 32'b11001101100110101101110101100100;
		#400 //-60957.91 * 0.00018769271 = -324775040.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110011101101100011110000001001;
		b = 32'b01001011101100010011100100101111;
		correct = 32'b00100111100000111001111010001011;
		#400 //8.485956e-08 * 23229022.0 = 3.6531697e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101101010010011000100110011000;
		b = 32'b00111010100000000000001100111010;
		correct = 32'b10110010010010011000010010000100;
		#400 //-1.1456079e-11 * 0.0009766587 = -1.172987e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100110111010001001110110101100;
		b = 32'b01001111111110101010110101001110;
		correct = 32'b01010110011011011000111000110000;
		#400 //5.4924878e+23 * 8411323400.0 = 65298737000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001111011011110111011111111111;
		b = 32'b00111110100101011011110010010011;
		correct = 32'b00010000010011001011010011000011;
		#400 //1.180672e-29 * 0.29245433 = 4.037116e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001100100101110000000010001110;
		b = 32'b00111001111110100101011000000110;
		correct = 32'b00010010000110100110101100101101;
		#400 //2.3265568e-31 * 0.00047747808 = 4.8725936e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100100101101101011011010111001;
		b = 32'b00111001001101000011100110010000;
		correct = 32'b00101011000000011100010010000111;
		#400 //7.923946e-17 * 0.00017187581 = 4.6102743e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111110000110011010101000110010;
		b = 32'b11010111001101001011110110110111;
		correct = 32'b11100110010110011010011001000010;
		#400 //5.1063897e+37 * -198726910000000.0 = -2.5695511e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010010001011000110001101110000;
		b = 32'b10000011111101011010111000101000;
		correct = 32'b11001101101100111010000100101001;
		#400 //5.4396196e-28 * -1.443979e-36 = -376710430.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011100100000101000100011110011;
		b = 32'b01011011000001110011010001010011;
		correct = 32'b00000000111101110010100010100100;
		#400 //8.638079e-22 * 3.8056653e+16 = 2.2697947e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111111110010111010100100101101;
		b = 32'b10111010000110010001110010010100;
		correct = 32'b11111111110010111010100100101101;
		#400 //nan * -0.0005840745 = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100101001011001001010000111011;
		b = 32'b10111110110000101100110101101111;
		correct = 32'b11100101111000101100101110000110;
		#400 //5.093634e+22 * -0.38047358 = -1.3387615e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011100010101010011000111001100;
		b = 32'b10000011111100010111011100001011;
		correct = 32'b11010111111000100000011100011100;
		#400 //7.054015e-22 * -1.4192038e-36 = -497040320000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010001011010101010000111100001;
		b = 32'b11000110100011011101100110101100;
		correct = 32'b01001010010100111011100100001010;
		#400 //-62983640000.0 * -18156.836 = 3468866.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000011000101110010010011011001;
		b = 32'b10001001011001010010001100000011;
		correct = 32'b11111001001010001101110100010010;
		#400 //151.14394 * -2.7581335e-33 = -5.4799357e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000001110010001010110111101111;
		b = 32'b10110001010000100101101001000100;
		correct = 32'b01010000000001000010101010110101;
		#400 //-25.084929 * -2.8282026e-09 = 8869565000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101110000010011101010000011001;
		b = 32'b01001100100011011011010101100000;
		correct = 32'b00100000111110001111110110011111;
		#400 //3.1338574e-11 * 74296060.0 = 4.2180667e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001100101011110010010010001100;
		b = 32'b10101011010000010101111100010001;
		correct = 32'b01100000111001111101111000011001;
		#400 //-91825250.0 * -6.8699305e-13 = 1.3366255e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011111001001010111100010011010;
		b = 32'b10110000001010100110011110110101;
		correct = 32'b01101110011110001001011001101111;
		#400 //-1.1923449e+19 * -6.1993016e-10 = 1.9233536e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101101110010101001001001000001;
		b = 32'b10110101100000011110000001001011;
		correct = 32'b01110111110001111010010100100001;
		#400 //-7.836598e+27 * -9.676527e-07 = 8.098565e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100110110101001101111111000100;
		b = 32'b00100101111111010000010011100101;
		correct = 32'b11000000010101110110000111001011;
		#400 //-1.4771107e-15 * 4.389182e-16 = -3.3653438
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101111110110100111001011000001;
		b = 32'b10001100011111111010111110101101;
		correct = 32'b01100010110110101011011101100001;
		#400 //-3.9735507e-10 * -1.9697351e-31 = 2.017302e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100000011111000010010111000110;
		b = 32'b00001011010001110101111111000100;
		correct = 32'b11010100101000011110000110001101;
		#400 //-2.1357728e-19 * 3.8398052e-32 = -5562191000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100000110001001010000101010110;
		b = 32'b11000111110010000110010011001101;
		correct = 32'b10011000011110110011000100110000;
		#400 //3.3310455e-19 * -102601.6 = -3.2465823e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001111100111111110001001111100;
		b = 32'b11100010100000110011001100001100;
		correct = 32'b00101100100110111111110001011101;
		#400 //-5364840400.0 * -1.2101009e+21 = 4.433383e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011001001110111001010011000011;
		b = 32'b01000111101101010010001101011111;
		correct = 32'b10010001000001001000110110001000;
		#400 //-9.6977156e-24 * 92742.74 = -1.0456577e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000010100101001001111111100100;
		b = 32'b11110111101101101110101100101011;
		correct = 32'b10001010010100000000000100100101;
		#400 //74.31229 * -7.420061e+33 = -1.0015051e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111001001110110101011100010;
		b = 32'b11110001100010011100100010011011;
		correct = 32'b00000101000110111000011110011001;
		#400 //-9.978861e-06 * -1.3645428e+30 = 7.31297e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001101010100101010110010010001;
		b = 32'b10111010111100001111010100010000;
		correct = 32'b11010001110111111101001110000110;
		#400 //220907790.0 * -0.0018383581 = -120165810000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011001101100111001011101011001;
		b = 32'b10011111000110000000010010010100;
		correct = 32'b01111010000101110011011110000111;
		#400 //-6318803700000000.0 * -3.219104e-20 = 1.9629076e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110100010100110010100011001111;
		b = 32'b11011101000101011011001001011001;
		correct = 32'b10010110101101001000110111110010;
		#400 //1.9665752e-07 * -6.741739e+17 = -2.9170148e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010001100111111010101001101;
		b = 32'b01101110100100010001001000100010;
		correct = 32'b10001011000111101100100000110111;
		#400 //-0.0006864861 * 2.2448624e+28 = -3.0580318e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010101011001000101010101000101;
		b = 32'b10010100111000110001101010010101;
		correct = 32'b11000000000000001011000101011101;
		#400 //4.61115e-26 * -2.2931627e-26 = -2.0108254
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100101000100100000000110100010;
		b = 32'b11000000111111010011110010000101;
		correct = 32'b00100011100100111001100110001010;
		#400 //-1.2664035e-16 * -7.9136376 = 1.6002798e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011111111111101001010011010000;
		b = 32'b11010010000000111111111001001101;
		correct = 32'b01001101011101101110000100001111;
		#400 //-3.6689032e+19 * -141726800000.0 = 258871540.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101101111000110101100100110110;
		b = 32'b11011111000111100001110001100001;
		correct = 32'b01001110001110000000110101001010;
		#400 //-8.7951183e+27 * -1.1393088e+19 = 771969660.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101101010111010010110000110000;
		b = 32'b11100000010110000010001100011110;
		correct = 32'b11001100100000101111101101101001;
		#400 //4.2781004e+27 * -6.22973e+19 = -68672330.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110110000111101011000001011101;
		b = 32'b11101110001010000001110010101000;
		correct = 32'b10000111011100011010011010010011;
		#400 //2.3646492e-06 * -1.3007031e+28 = -1.8179777e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101100110100011101101000100111;
		b = 32'b11000010000101000000011111001101;
		correct = 32'b00101010001101010111010011010110;
		#400 //-5.964357e-12 * -37.007618 = 1.6116565e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010101110000110111101011001001;
		b = 32'b11111110100000111010110110100011;
		correct = 32'b10010110101111100000010011100111;
		#400 //26866516000000.0 * -8.751522e+37 = -3.069925e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011010010100100100010000110001;
		b = 32'b01001110111111111000001101100101;
		correct = 32'b11001010110100101010101010111011;
		#400 //-1.4796181e+16 * 2143400600.0 = -6903133.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011111001100100111001101010001;
		b = 32'b01111111110011110111010001111110;
		correct = 32'b01111111110011110111010001111110;
		#400 //3.7788354e-20 * nan = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000110011000001001011111001110;
		b = 32'b01001000100001000011001011000110;
		correct = 32'b00111101010110010111010111011101;
		#400 //14373.951 * 270742.2 = 0.05309092
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011111110101001001110011101001;
		b = 32'b11111111110111010100011001011001;
		correct = 32'b11111111110111010100011001011001;
		#400 //-3.0640752e+19 * nan = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000010011110100010011110101001;
		b = 32'b11110011000001101000110001100010;
		correct = 32'b00001110111011011111101011100110;
		#400 //-62.53873 * -1.066002e+31 = 5.8666617e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110110011100100011011110111010;
		b = 32'b11011101000001110100001000111100;
		correct = 32'b01011000111001010011100000001101;
		#400 //-1.22818956e+33 * -6.0915116e+17 = 2016231200000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000010110011110000011100001101;
		b = 32'b11110110100111010101111000100010;
		correct = 32'b00001011101010000110010001110100;
		#400 //-103.51377 * -1.5958981e+33 = 6.486239e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111011101101111111100000100000;
		b = 32'b11000101110101010111010101110110;
		correct = 32'b11110101010111001010001000011111;
		#400 //1.9104458e+36 * -6830.6826 = -2.7968592e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101010100001011001101010011110;
		b = 32'b00011100100010011101101011010001;
		correct = 32'b01001101011110000001101100101111;
		#400 //2.3732833e-13 * 9.122462e-22 = 260158190.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010001001011001011111001010101;
		b = 32'b11001010010000111011100001110111;
		correct = 32'b10000110011000011111001000111111;
		#400 //1.3627058e-28 * -3206685.8 = -4.249577e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100010010010011001111001001010;
		b = 32'b10011111110110010101110100110100;
		correct = 32'b01000001111011010111010010011010;
		#400 //-2.7324377e-18 * -9.2057266e-20 = 29.681934
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010000001101001100101110011101;
		b = 32'b00011100010100100110101111000000;
		correct = 32'b00110011010110111111010100010010;
		#400 //3.56556e-29 * 6.9622435e-22 = 5.12128e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110100101011001000110000011000;
		b = 32'b01101110110000011111000011110111;
		correct = 32'b01000101011000111100001010011010;
		#400 //1.0936481e+32 * 3.0010958e+28 = 3644.1626
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010011011001001101011000001011;
		b = 32'b11110110010110111110101001011011;
		correct = 32'b10011100100001010011000100110100;
		#400 //982843600000.0 * -1.1151038e+33 = -8.81392e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111010011110011101000100000000;
		b = 32'b01001010100001100000111011000100;
		correct = 32'b11101111011011101000011100100110;
		#400 //-3.2428024e+35 * 4392802.0 = -7.3820817e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010110010111010011101101011100;
		b = 32'b10100010011010100010100001010000;
		correct = 32'b00110011011100011101111001100010;
		#400 //-1.7870968e-25 * -3.1734255e-18 = 5.631444e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001001100110001101110101000100;
		b = 32'b11011001000000111110101000000000;
		correct = 32'b10110000000101000101010000100001;
		#400 //1252264.5 * -2320656700000000.0 = -5.396164e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111101100110001010100111010101;
		b = 32'b01100111100000111101000110111101;
		correct = 32'b00010101100101000011110101111101;
		#400 //0.07454268 * 1.244998e+24 = 5.9873735e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100100010111000110111011001;
		b = 32'b10010011101001011111100000111001;
		correct = 32'b11110000010101110100000101011110;
		#400 //1116.4327 * -4.1896622e-27 = -2.664732e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100001011110101011110110101000;
		b = 32'b00001111011111100010101011010111;
		correct = 32'b11010001011111001000110001111110;
		#400 //-8.4954303e-19 * 1.25314175e-29 = -67793050000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110010001101010010100110011100;
		b = 32'b01110111111001100000111110111010;
		correct = 32'b00111001110010011001011010000011;
		#400 //3.5882937e+30 * 9.3324004e+33 = 0.00038449847
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110001101111001101101110101100;
		b = 32'b10001101000100110001100000101010;
		correct = 32'b11100100001001000101011110100011;
		#400 //5.496494e-09 * -4.532696e-31 = -1.2126324e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100111101100110010001011001010;
		b = 32'b00110101100110011001011111111101;
		correct = 32'b10110001100101010100100100111001;
		#400 //-4.97202e-15 * 1.1443623e-06 = -4.344795e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110000001001100111000101011100;
		b = 32'b10110001100100000110100110001100;
		correct = 32'b10111110000100111000011011011011;
		#400 //6.055154e-10 * -4.202951e-09 = -0.14406912
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001011010101100010111110110101;
		b = 32'b01000111000010111010111111001101;
		correct = 32'b00000011110001000100010001000111;
		#400 //4.1250792e-32 * 35759.8 = 1.153552e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010011101111010000010110010110;
		b = 32'b10010011010111011100001000111011;
		correct = 32'b10111111110110100011010101010001;
		#400 //4.7715816e-27 * -2.7989885e-27 = -1.7047521
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101010000111110010010111110110;
		b = 32'b00110100111010110111010010111000;
		correct = 32'b10110100101011010000100011001010;
		#400 //-1.4135207e-13 * 4.3857085e-07 = -3.2230156e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000110100111000011111000001000;
		b = 32'b01110101101100101111101100010110;
		correct = 32'b00010000010111110111101000000110;
		#400 //19999.016 * 4.5377025e+32 = 4.4073e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010010010111100111101000010101;
		b = 32'b01111010000110011110000101001010;
		correct = 32'b00010111101110010000111101011101;
		#400 //238882730000.0 * 1.997477e+35 = 1.1959223e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110011011101000100111110011101;
		b = 32'b00001011000010000101010100000001;
		correct = 32'b11100111111001010110000100110101;
		#400 //-5.6883085e-08 * 2.6256597e-32 = -2.1664302e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011110001011100100111011010;
		b = 32'b10110111011110010011000100101101;
		correct = 32'b01010011110010110011000100101010;
		#400 //-25924532.0 * -1.4853006e-05 = 1745406400000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101001100011001010100111100111;
		b = 32'b11110111011000011000110000000110;
		correct = 32'b10110001100111111010011111101001;
		#400 //2.1256494e+25 * -4.574636e+33 = -4.646598e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011110001011111001000100110000;
		b = 32'b10111101110011011110110011000111;
		correct = 32'b01011111110110100100001010010101;
		#400 //-3.1627364e+18 * -0.10054927 = 3.1454593e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010100110111110011001111100101;
		b = 32'b10010101110101001111110101110000;
		correct = 32'b00111110100001100010001100110100;
		#400 //-2.2537714e-26 * -8.602597e-26 = 0.26198733
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100000101011000100101011010001;
		b = 32'b00011101010011110010000111001000;
		correct = 32'b01000010110101001111000011001111;
		#400 //2.9187443e-19 * 2.7413686e-21 = 106.47033
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110100011010111100101010011110;
		b = 32'b11110001111000011110100010101001;
		correct = 32'b10000010000001011001100101111001;
		#400 //2.1959792e-07 * -2.2372927e+30 = -9.815341e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111011011111011001101101000101;
		b = 32'b01101000011110100101010110100110;
		correct = 32'b01010010100000011010110001001010;
		#400 //1.31680035e+36 * 4.7286862e+24 = 278470660000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100110000110010011010010101100;
		b = 32'b01010100000001010101010010010000;
		correct = 32'b00010001100100110001010010110010;
		#400 //5.315392e-16 * 2290597500000.0 = 2.3205265e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010111111000111001011010000110;
		b = 32'b11000101101110011010111101010000;
		correct = 32'b01010001100111001110001010110011;
		#400 //-500471270000000.0 * -5941.914 = 84227285000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111100110010000101100101100001;
		b = 32'b01011101000010110010001011110101;
		correct = 32'b11011111001110000101000000101000;
		#400 //-8.3221775e+36 * 6.266153e+17 = -1.3281159e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001111100000011001001000111110;
		b = 32'b10101010001111101000100111001010;
		correct = 32'b10100100101011100001011001001010;
		#400 //1.2776713e-29 * -1.6923195e-13 = -7.549823e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100001010001010111110100011011;
		b = 32'b00101001000101011100000111110010;
		correct = 32'b10110111101010001100101111100101;
		#400 //-6.691177e-19 * 3.3252867e-14 = -2.0122106e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101101010101111110110100111001;
		b = 32'b10111110000010101010110110011001;
		correct = 32'b10101110110001110100110011101010;
		#400 //1.2274009e-11 * -0.13542785 = -9.063135e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000010101011110010011010101111;
		b = 32'b00010011100110110010001001001101;
		correct = 32'b01101110100100001000010000011000;
		#400 //87.575554 * 3.9161324e-27 = 2.2362766e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000011101111001010110111101010;
		b = 32'b10001010001011100010010111000001;
		correct = 32'b11111001000010101010111001011010;
		#400 //377.3587 * -8.384896e-33 = -4.5004577e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111011010010000000010001100111;
		b = 32'b11000111100100100001111111111011;
		correct = 32'b01110011001011110011010100100111;
		#400 //-1.0385487e+36 * -74815.96 = 1.3881378e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101111101100010001111110001100;
		b = 32'b00101010001101010110101001011100;
		correct = 32'b11000100111110011111000101110000;
		#400 //-3.2218528e-10 * 1.611293e-13 = -1999.5449
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011111000101011010000101110000;
		b = 32'b01111110110011100000010110111000;
		correct = 32'b00011111101110011110110110110110;
		#400 //1.0782022e+19 * 1.3692533e+38 = 7.874381e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001110010110010110110101010101;
		b = 32'b00001111101010111001111100101001;
		correct = 32'b11111110001000100010100110110000;
		#400 //-911955260.0 * 1.6923208e-29 = -5.3887847e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001110101001101101010101001010;
		b = 32'b10011111001111110000110111011010;
		correct = 32'b11101110110111111000101110100111;
		#400 //1399498000.0 * -4.045728e-20 = -3.4591993e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010101001001010110000100010010;
		b = 32'b01010000110101110001111000110100;
		correct = 32'b00000011110001001100111100000001;
		#400 //3.339806e-26 * 28872647000.0 = 1.156737e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001111101110100011010001101010;
		b = 32'b10100001000010101111100010010101;
		correct = 32'b01101110001010111000000100111111;
		#400 //-6247994400.0 * -4.7085214e-19 = 1.3269546e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000110100110110001011101110111;
		b = 32'b00010110001100011010001010001100;
		correct = 32'b01101111110111111000001011110110;
		#400 //19851.732 * 1.4349237e-25 = 1.3834696e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111100110010011010000001111001;
		b = 32'b01110110111001100010001100110100;
		correct = 32'b00000101011000000100100100001101;
		#400 //0.024612652 * 2.3338716e+33 = 1.0545847e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000011011111110000100100011000;
		b = 32'b01000100101011000001111010001001;
		correct = 32'b00111110001111011010100110010000;
		#400 //255.03552 * 1376.9542 = 0.18521714
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000001101101101100011000101101;
		b = 32'b10000111110011010000010001100010;
		correct = 32'b11111001011001000011100111000111;
		#400 //22.846766 * -3.0847548e-34 = -7.406347e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100101010001010010110110110001;
		b = 32'b10101001100110000000010111011000;
		correct = 32'b01111011001001100000010100100110;
		#400 //-5.8196816e+22 * -6.75117e-14 = 8.620257e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100011001000101000101100111111;
		b = 32'b11011000000010100110101001100000;
		correct = 32'b01001010100101100101000000010011;
		#400 //-2.9984063e+21 * -608757900000000.0 = 4925449.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110011010001011001000000010011;
		b = 32'b10110100010011101101111101101101;
		correct = 32'b11111110011101000111101010101001;
		#400 //1.5652537e+31 * -1.9266527e-07 = -8.124213e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011100100111010101001110001100;
		b = 32'b01111011111000001101000101111001;
		correct = 32'b00100000001100110010010110101011;
		#400 //3.5426746e+17 * 2.3346462e+36 = 1.5174353e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001101000100110001001100000101;
		b = 32'b01001000000010101000010101011001;
		correct = 32'b11000100100001111110011101011101;
		#400 //-154218580.0 * 141845.39 = -1087.2301
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011101100101011101111101100110;
		b = 32'b00011110011101101100010011100011;
		correct = 32'b00111110100110110111101010011100;
		#400 //3.967096e-21 * 1.3063847e-20 = 0.3036698
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001110010000101101000000111111;
		b = 32'b01010101011100001101110011100010;
		correct = 32'b00111000010011110000111010000000;
		#400 //817106900.0 * 16551967000000.0 = 4.936615e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101101010001011011101000101111;
		b = 32'b01000100100111110000110001001001;
		correct = 32'b00101000000111110010000011101111;
		#400 //1.1239495e-11 * 1272.3839 = 8.833414e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001001000100011111101101100111;
		b = 32'b00101001000111001100010000010110;
		correct = 32'b10011111011011100110001111001000;
		#400 //-1.7571949e-33 * 3.4809036e-14 = -5.0480997e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001100110101000011000111100101;
		b = 32'b10111011100000111011001110000101;
		correct = 32'b10010000110011100011101101000100;
		#400 //3.26938e-31 * -0.004019203 = -8.1343986e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110100010111010100011100111001;
		b = 32'b01110010001000100000000000000111;
		correct = 32'b01000001101011101101011001000101;
		#400 //7.0125865e+31 * 3.2087427e+30 = 21.854624
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111111010000000100110011100001;
		b = 32'b01111111010101000001000100001100;
		correct = 32'b10111111011010000010001110000111;
		#400 //-2.5561095e+38 * 2.8188485e+38 = -0.9067921
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010000101001000010110110001110;
		b = 32'b10100000111001110011100111100111;
		correct = 32'b11101111001101011100010010100101;
		#400 //22035591000.0 * -3.917124e-19 = -5.6254515e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101111001010010011010000011001;
		b = 32'b10110000110111011001100101001010;
		correct = 32'b10111101110000110111100010001000;
		#400 //1.5388969e-10 * -1.6123434e-09 = -0.09544474
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100001010010100100000011000111;
		b = 32'b00100100010110110100110111110000;
		correct = 32'b00111100011011000001100001101110;
		#400 //6.8525994e-19 * 4.755407e-17 = 0.014410121
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101110111000001111010001011111;
		b = 32'b01110110111001100110001010111111;
		correct = 32'b00110111011110011111011100001011;
		#400 //3.4810034e+28 * 2.3363888e+33 = 1.4899076e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101001000010101110100011110010;
		b = 32'b01100100100001100000101100010000;
		correct = 32'b01000100000001001010010110110111;
		#400 //1.0495739e+25 * 1.9781287e+22 = 530.5893
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111101100110101110100110000010;
		b = 32'b00011010100010000011010001111111;
		correct = 32'b11100010100100011001010010000101;
		#400 //-0.07564069 * 5.6333094e-23 = -1.3427399e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010101110101011110100000100101;
		b = 32'b00010001000000010100111101111010;
		correct = 32'b01000100010100111011110100110010;
		#400 //8.6396274e-26 * 1.0200796e-28 = 846.9562
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110000111101001111001000100100;
		b = 32'b01111001010000101110001100101110;
		correct = 32'b00110111001000001110000010111011;
		#400 //6.0645658e+29 * 6.3244584e+34 = 9.589067e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011101001010001000100000101000;
		b = 32'b01111101101001001001101111010100;
		correct = 32'b00011111000000110000110011111000;
		#400 //7.59e+17 * 2.7350312e+37 = 2.7751057e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111100010010011001111001001001;
		b = 32'b10100001100010000100111111111111;
		correct = 32'b11011010001111010101001011001010;
		#400 //0.0123058045 * -9.236893e-19 = -1.332245e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111001010011110100101001110;
		b = 32'b11001011010001100111100100001011;
		correct = 32'b00101011010110110010100011110110;
		#400 //-1.0127505e-05 * -13007115.0 = 7.7861274e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101110101010001000001101010101;
		b = 32'b10011101100111101110110011001010;
		correct = 32'b11010000100001111011100011101011;
		#400 //7.663085e-11 * -4.2067086e-21 = -18216344000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110101011000101010111010101100;
		b = 32'b00111110110010110110111010010011;
		correct = 32'b00110110000011101010000100010100;
		#400 //8.444574e-07 * 0.397328 = 2.1253409e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001000110110000000101111101010;
		b = 32'b10001010111000010100101000011001;
		correct = 32'b00111101011101010111111101000101;
		#400 //-1.3002828e-33 * -2.1694584e-32 = 0.059935827
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111010011010001101000011010110;
		b = 32'b01111101100011101011100100000010;
		correct = 32'b00111100010100001100110010101001;
		#400 //3.0221214e+35 * 2.3713874e+37 = 0.012744107
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110010100101100100100001001111;
		b = 32'b01010100011100011111011100111010;
		correct = 32'b00011101100111101111111110111110;
		#400 //1.749518e-08 * 4156939600000.0 = 4.2086683e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011000101001111101000001011001;
		b = 32'b00100110000001011011101011110110;
		correct = 32'b01110010001000001001111110000001;
		#400 //1476106300000000.0 * 4.6397024e-16 = 3.1814675e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111011110111001000011001100001;
		b = 32'b11101111000001111100101111010010;
		correct = 32'b11001100010011111101110101001001;
		#400 //2.2900617e+36 * -4.202688e+28 = -54490404.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011100101011010110011010001101;
		b = 32'b00001010110000110110100001010110;
		correct = 32'b11010001011000110010101101000111;
		#400 //-1.1474688e-21 * 1.8817064e-32 = -60980230000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110010000010000011111101001100;
		b = 32'b11001100100001111101101011000111;
		correct = 32'b00100101000000000101111010110101;
		#400 //-7.930634e-09 * -71226936.0 = 1.1134318e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110000000111100011110001101000;
		b = 32'b01000101101001100010111110001101;
		correct = 32'b00101001111100111100000011111001;
		#400 //5.756591e-10 * 5317.944 = 1.0824843e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111101101110011000101000110101;
		b = 32'b01000101110000000000101101110010;
		correct = 32'b00110111011101110101010000110011;
		#400 //0.09059564 * 6145.4307 = 1.4741951e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001001001110011100010010111000;
		b = 32'b10001111001110011011011100110010;
		correct = 32'b01111001100000000000100101010010;
		#400 //-760907.5 * -9.156486e-30 = 8.310038e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001101011111011101000110111010;
		b = 32'b01001001000010100011000100010111;
		correct = 32'b00000011111010110001100110010001;
		#400 //7.8214093e-31 * 566033.44 = 1.3817928e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111000101010000100110101001;
		b = 32'b11101111010010001101010010001110;
		correct = 32'b10010111001111011111101011001000;
		#400 //38153.66 * -6.2153965e+28 = -6.1385724e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010100111001011011101101000100;
		b = 32'b00111011001111011101001000101001;
		correct = 32'b10011001000110101110100110011000;
		#400 //-2.3196954e-26 * 0.0028964377 = -8.008787e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000011011111001111010110000000;
		b = 32'b00011111010101010000010101000111;
		correct = 32'b10100011100101111111111110001010;
		#400 //-7.4337964e-37 * 4.510887e-20 = -1.6479678e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101101001001110011111000010011;
		b = 32'b11010010111110111001000110001000;
		correct = 32'b01011001101010100011000001000101;
		#400 //-3.23494e+27 * -540239200000.0 = 5987977400000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000001110011100001000010110111;
		b = 32'b10000101010110010101001001010110;
		correct = 32'b00111011111100101011110110000100;
		#400 //-7.5696433e-38 * -1.0218414e-35 = 0.007407846
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100011010111101011100100000100;
		b = 32'b11000000000111101010101110101100;
		correct = 32'b10100010101100111010101111001000;
		#400 //1.2073823e-17 * -2.479228 = -4.8699928e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000111101010000000101100010011;
		b = 32'b00011111100001011011111111110001;
		correct = 32'b00100111101000001101000110111010;
		#400 //2.528434e-34 * 5.664523e-20 = 4.4636307e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001110100100001110010100001011;
		b = 32'b10010100001010110100100111001010;
		correct = 32'b10111001110110001000110110101001;
		#400 //3.57193e-30 * -8.647846e-27 = -0.00041304276
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010110010000100010010001101010;
		b = 32'b10001001100111001010111110011011;
		correct = 32'b11001100000111101001100101001100;
		#400 //1.5682685e-25 * -3.7720773e-33 = -41575730.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010100110010101010001001100011;
		b = 32'b11111100101101001101110001100110;
		correct = 32'b00010111100011110110100011011011;
		#400 //-6962462300000.0 * -7.512669e+36 = 9.267628e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010001000111101000110110010011;
		b = 32'b11110111101011101000101001101011;
		correct = 32'b10011000111010001000110100000000;
		#400 //42561253000.0 * -7.080212e+33 = -6.0112968e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011100110111011100111100000001;
		b = 32'b11000001100011000010001100111000;
		correct = 32'b01011010110010101001100011101100;
		#400 //-4.994686e+17 * -17.517197 = 2.8513042e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000001011000110001010111000101;
		b = 32'b00111111010001100011001110110000;
		correct = 32'b10000001100100101010011100100101;
		#400 //-4.1708934e-38 * 0.7742262 = -5.387177e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111101010010101110000100111111;
		b = 32'b00110110110001111100001110010110;
		correct = 32'b11000110000000011111111100011011;
		#400 //-0.049531218 * 5.9534314e-06 = -8319.776
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010000000010001100001110011011;
		b = 32'b10111110010110101100011111000100;
		correct = 32'b00010001001000000000011111100111;
		#400 //-2.697196e-29 * -0.21365267 = 1.262421e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110110111010000110100000110110;
		b = 32'b01111101101110100000100111001010;
		correct = 32'b10111000100111111110011100110111;
		#400 //-2.3568877e+33 * 3.0910904e+37 = -7.624778e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011111100100101010100100001010;
		b = 32'b10100000100100110010001111010110;
		correct = 32'b11111110011111110010101001011010;
		#400 //2.1135978e+19 * -2.4926483e-19 = -8.479326e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011011101111100000001100001010;
		b = 32'b00101001010100110001000101111000;
		correct = 32'b01110001111001100111011000010001;
		#400 //1.0696717e+17 * 4.6866563e-14 = 2.2823771e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100110000010001001100101110001;
		b = 32'b10000010100111011100001000101111;
		correct = 32'b11100010110111011010101000010011;
		#400 //4.739243e-16 * -2.3180533e-37 = -2.0444928e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010111000111110110010110011100;
		b = 32'b10010101011110101011000100110001;
		correct = 32'b11000001001000101100010110010100;
		#400 //5.150392e-25 * -5.0626877e-26 = -10.173237
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101101000000110111000011000010;
		b = 32'b01101000111001010000101000001111;
		correct = 32'b11000011100100101110100110100000;
		#400 //-2.5424283e+27 * 8.65286e+24 = -293.8252
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101010101101100000111110110100;
		b = 32'b01000010000111011010100100000000;
		correct = 32'b00101000000100111100111110000111;
		#400 //3.234059e-13 * 39.41504 = 8.2051396e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101101011110001101100000011110;
		b = 32'b10011111010000100011100100110111;
		correct = 32'b01001101101000111111111100110111;
		#400 //-1.41451555e-11 * -4.1128425e-20 = 343926500.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111011100111001010001111011;
		b = 32'b00111111010011101000101100111111;
		correct = 32'b10110111100101101111001110111101;
		#400 //-1.45184995e-05 * 0.8068122 = -1.7994893e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100111100110001100001110110;
		b = 32'b01011001011101111101000111101111;
		correct = 32'b00101010111110110001111010011011;
		#400 //1944.7644 * 4359696500000000.0 = 4.4607793e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101010101001010001011011011000;
		b = 32'b00100101110101101100101011011110;
		correct = 32'b01000100010001001100001011100101;
		#400 //2.932574e-13 * 3.726055e-16 = 787.0452
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011000101001111110100101000011;
		b = 32'b10110111000101101111011110101110;
		correct = 32'b00100001000011100101110110101111;
		#400 //-4.3404022e-24 * -8.998364e-06 = 4.823546e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001001110010100101101000011110;
		b = 32'b00011101100101110100101111001110;
		correct = 32'b11101011101010110011000111001001;
		#400 //-1657667.8 * 4.0047747e-21 = -4.1392284e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110010000001001010111100011;
		b = 32'b11101000000001000010111001110111;
		correct = 32'b10010101101110100111111000111110;
		#400 //0.18807177 * -2.496838e+24 = -7.5323977e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001011010100001011010101111001;
		b = 32'b11001001001000111001101011101100;
		correct = 32'b00000001101000110100100110110001;
		#400 //-4.0195868e-32 * -670126.75 = 5.9982485e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100001011110100100010100100000;
		b = 32'b11001100001111001000010001110101;
		correct = 32'b00010100101010011110110111001111;
		#400 //-8.479478e-19 * -49418708.0 = 1.7158438e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011001011001010110100101011110;
		b = 32'b11001001000011010000111110101100;
		correct = 32'b11001111110100000010101101110111;
		#400 //4035851400000000.0 * -577786.75 = -6985019000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101010011011110100100001111001;
		b = 32'b10111010001001011100011001111110;
		correct = 32'b10101111101110001100000111101010;
		#400 //2.1252608e-13 * -0.0006323828 = -3.360719e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010000010100011000001011100000;
		b = 32'b11001110011111001110001001100110;
		correct = 32'b11000001010101000001011110101101;
		#400 //14060061000.0 * -1060673900.0 = -13.25578
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000101001011101100101101000100;
		b = 32'b00001111011001000001101011101101;
		correct = 32'b11110101010001000010101101100001;
		#400 //-2796.704 * 1.12464536e-29 = -2.4867432e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110000000101100011101001110011;
		b = 32'b10111011010101101110010110010111;
		correct = 32'b01110100001100101111011001011111;
		#400 //-1.8597365e+29 * -0.0032790655 = 5.6715444e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000010001111001001010010010000;
		b = 32'b11011100010111111111010110011111;
		correct = 32'b10100101010101111000111100110100;
		#400 //47.14508 * -2.5215593e+17 = -1.8696796e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011101011110000010111101000011;
		b = 32'b00001111001011000000000010101011;
		correct = 32'b11001101101110001011000101010111;
		#400 //-3.284696e-21 * 8.4803834e-30 = -387328740.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000101100010000111111010100100;
		b = 32'b01000101100111000111000100100010;
		correct = 32'b00111111010111110101101111001010;
		#400 //4367.83 * 5006.1416 = 0.87249434
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101110100101000111000010011100;
		b = 32'b01010110101001011110100001001011;
		correct = 32'b11010111011001010000110000001111;
		#400 //-2.296996e+28 * 91208555000000.0 = -251839950000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000010011111001100011001111101;
		b = 32'b01110011010010000101001010101111;
		correct = 32'b00001110101000011000001111110000;
		#400 //63.193836 * 1.5871222e+31 = 3.9816615e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011011001110101111101001010110;
		b = 32'b00110100100001011001011101110001;
		correct = 32'b10100110001100110010011011011011;
		#400 //-1.5466447e-22 * 2.488337e-07 = -6.215576e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011001101000100111101001100;
		b = 32'b10011111001000010110011110101110;
		correct = 32'b01101011100011101111110111111110;
		#400 //-11816780.0 * -3.4178838e-20 = 3.4573382e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010100101100010111101000000100;
		b = 32'b00111001000001001101001110111100;
		correct = 32'b10011011001010110000011011100100;
		#400 //-1.792056e-26 * 0.00012667378 = -1.4147015e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101100011101010110000011110111;
		b = 32'b01011010001101101110000001110001;
		correct = 32'b10010001101010111011111100101011;
		#400 //-3.487042e-12 * 1.2868805e+16 = -2.709686e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011100111101111111111001101110;
		b = 32'b11001010111100110000001011110001;
		correct = 32'b01010001100000101001111111010101;
		#400 //-5.5843254e+17 * -7963000.5 = 70128410000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010111010001000000100111000101;
		b = 32'b00011010101001001001000101000000;
		correct = 32'b11111100000110000111101001010110;
		#400 //-215546240000000.0 * 6.8063474e-23 = -3.1668416e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001000000100111011011110010001;
		b = 32'b10001010100100101101001101000011;
		correct = 32'b10111101000000001100011100001000;
		#400 //4.4451985e-34 * -1.4138756e-32 = -0.03143981
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110100000011010101111001100001;
		b = 32'b11001100010001110110000001100010;
		correct = 32'b01100111001101011000010010001101;
		#400 //-4.480152e+31 * -52265350.0 = 8.5719346e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010001101011100110001110000100;
		b = 32'b00111010111111101010000101111011;
		correct = 32'b11010110001011110101001110010011;
		#400 //-93624240000.0 * 0.0019426787 = -48193370000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100111111011001011110101111;
		b = 32'b10101101100001001011010101100100;
		correct = 32'b11010110111101001001100001001110;
		#400 //2028.7401 * -1.5087216e-11 = -134467490000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100010110101110011001100100111;
		b = 32'b10000010100001111111111111000111;
		correct = 32'b11011111110010101000101011010100;
		#400 //5.8330026e-18 * -1.9983276e-37 = -2.9189421e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010001111100011101110011001110;
		b = 32'b11101100100011001000110010101000;
		correct = 32'b10100100110111000100010001011010;
		#400 //129848950000.0 * -1.3593108e+27 = -9.552558e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111011101111100010110011100000;
		b = 32'b00111111110111100111011100001001;
		correct = 32'b01111011010110101101011111000110;
		#400 //1.9748932e+36 * 1.7380077 = 1.1362971e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011111000010110011010011000000;
		b = 32'b11111001110001000000000000010111;
		correct = 32'b00100100101101011101000111100000;
		#400 //-1.0030853e+19 * -1.272115e+35 = 7.885178e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001101000111110000111011100001;
		b = 32'b10010100100101010110111111100111;
		correct = 32'b10111000000010000011110110101000;
		#400 //4.9013568e-31 * -1.5089293e-26 = -3.248235e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000110001101000011101000001100;
		b = 32'b01111111110011101101000000111111;
		correct = 32'b01111111110011101101000000111111;
		#400 //-11534.512 * nan = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000000011000000001011111011101;
		b = 32'b00110011010000111110010011001011;
		correct = 32'b00001100011110110010011110111011;
		#400 //8.824768e-39 * 4.561006e-08 = 1.9348293e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111000100100001110100101100101;
		b = 32'b11110111011000000010001010111101;
		correct = 32'b11000000101001011000001101011011;
		#400 //2.3513267e+34 * -4.546012e+33 = -5.1722846
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101001101100000100110100001001;
		b = 32'b01111011100011111101101101011100;
		correct = 32'b00101101100111001101111000101011;
		#400 //2.6641842e+25 * 1.4938952e+36 = 1.7833809e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110101011111011110110011000010;
		b = 32'b10000111001110011011101100100101;
		correct = 32'b11101101101011101111111100111101;
		#400 //9.459437e-07 * -1.397285e-34 = -6.7698695e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011000100011101000100111001001;
		b = 32'b11000011000001011101010110011100;
		correct = 32'b01010101000010000101001100001010;
		#400 //-1253779500000000.0 * -133.83441 = 9368139000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011110001100101011110001001101;
		b = 32'b11000101111010010101000101110011;
		correct = 32'b10010111110001000001110001110111;
		#400 //9.462181e-21 * -7466.181 = -1.2673389e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010001010101000001100001001101;
		b = 32'b11000010110000100110101101110011;
		correct = 32'b01001110000010111010001100000110;
		#400 //-56933798000.0 * -97.20986 = 585679200.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100001110110101101001000100001;
		b = 32'b11111101011111111011100111001101;
		correct = 32'b10100011110110110000111000110011;
		#400 //5.0456645e+20 * -2.1244867e+37 = -2.3750041e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000010110100010010010000000100;
		b = 32'b00110010111000001001011100110000;
		correct = 32'b01001111011011100110001110110001;
		#400 //104.57034 * 2.6145784e-08 = 3999510800.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101010000100000000100110011110;
		b = 32'b10011000000000000111100111100100;
		correct = 32'b11010001100011111000000011110110;
		#400 //1.2793106e-13 * -1.6605151e-24 = -77042990000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001000000100110010100101100100;
		b = 32'b11100101101010101111001010010011;
		correct = 32'b00100001110111000110000100111100;
		#400 //-150693.56 * -1.0090963e+23 = 1.4933518e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100000100001110111111001011001;
		b = 32'b11011101111111111010110010010001;
		correct = 32'b11000010000001111010101010010000;
		#400 //7.810671e+19 * -2.3029075e+18 = -33.916565
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110011000100000001111111101001;
		b = 32'b11100011010010001101000100101010;
		correct = 32'b10001111001101111011101010011110;
		#400 //3.3556635e-08 * -3.7044207e+21 = -9.058538e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011010000010011011010001110111;
		b = 32'b10011000010100100101110101000011;
		correct = 32'b01000001001001111001010000000011;
		#400 //-2.8476714e-23 * -2.7188949e-24 = 10.473636
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110011111110000010011001010000;
		b = 32'b10010011111001010010000101010110;
		correct = 32'b11011111100010101001111111111010;
		#400 //1.1555369e-07 * -5.78406e-27 = -1.9977955e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100100001001110011101010101001;
		b = 32'b11111001001010001110010010010011;
		correct = 32'b00101010011111010111101001101011;
		#400 //-1.2339333e+22 * -5.480887e+34 = 2.2513386e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101111011011111110100110001101;
		b = 32'b01100110100111110010001010000101;
		correct = 32'b11001000010000001111100100101010;
		#400 //-7.4249263e+28 * 3.7574652e+23 = -197604.66
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100111000101000101100000001010;
		b = 32'b01110100001010010100101100101010;
		correct = 32'b00110010011000000101001000010001;
		#400 //7.005343e+23 * 5.3651286e+31 = 1.3057176e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101101011110111001010001100011;
		b = 32'b11011010010000010111110110111001;
		correct = 32'b01010010101001100110110101100001;
		#400 //-4.866258e+27 * -1.3615726e+16 = 357399820000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010101100010000101111111111110;
		b = 32'b00110000010100010011100111000011;
		correct = 32'b11100100101001101101110011100110;
		#400 //-18743233000000.0 * 7.611584e-10 = -2.4624615e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100010010101001000101000010101;
		b = 32'b01000001110111000111000011110111;
		correct = 32'b11011111111101101101001011010000;
		#400 //-9.801649e+20 * 27.555159 = -3.5571013e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111001101001000000010010100001;
		b = 32'b10101100010000110110000010010101;
		correct = 32'b01001100110101101110100100010111;
		#400 //-0.00031283966 * -2.776478e-12 = 112675000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001100000001000001001001110111;
		b = 32'b11000100001101001001111101110011;
		correct = 32'b00000111001110110011000000101101;
		#400 //-1.0174467e-31 * -722.4914 = 1.4082474e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110000010101100111100001000110;
		b = 32'b10111010011011000010110001101110;
		correct = 32'b11110101011010000111100101101001;
		#400 //2.6550078e+29 * -0.0009009306 = -2.9469613e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101000010010010000110010011111;
		b = 32'b01011110010011101111011001100000;
		correct = 32'b01001001011110001010111110010100;
		#400 //3.797714e+24 * 3.7283032e+18 = 1018617.25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000001000000011101100011101001;
		b = 32'b11100111001000011110111000011101;
		correct = 32'b00011001010011010100011110000011;
		#400 //-8.115457 * -7.646934e+23 = 1.0612693e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101100111011001011000010111110;
		b = 32'b11010110100000000000000100011010;
		correct = 32'b11010101111011001010111010110101;
		#400 //2.2891291e+27 * -70371110000000.0 = -32529388000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110000011000110110110011000111;
		b = 32'b01100010010010100101000001001010;
		correct = 32'b00001101100011111110001100101111;
		#400 //8.27367e-10 * 9.330069e+20 = 8.867748e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000011001010010100101100100101;
		b = 32'b10011100010010001000010100010100;
		correct = 32'b01100110010110000010001001001011;
		#400 //-169.29353 * -6.634645e-22 = 2.5516594e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110100001100010010001010111100;
		b = 32'b00001000101110110100101100001100;
		correct = 32'b11101010111100100001110111001001;
		#400 //-1.6497046e-07 * 1.1272297e-33 = -1.4635035e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100101100100011111100101001111;
		b = 32'b10100011000101111101000100000101;
		correct = 32'b01000001111101100010010111011101;
		#400 //-2.5322428e-16 * -8.229988e-18 = 30.768488
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000101101100110111100100000010;
		b = 32'b00000101110110001001101000101101;
		correct = 32'b00111111010101000001110111110000;
		#400 //1.687753e-35 * 2.0369178e-35 = 0.8285818
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100001001010011110101111010100;
		b = 32'b01000110001111101111100111101001;
		correct = 32'b01011010011000111100011010110010;
		#400 //1.9590581e+20 * 12222.478 = 1.6028322e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011111110101101011100100011111;
		b = 32'b11001110110101110110111111100100;
		correct = 32'b10010000011111110010011011010001;
		#400 //9.093878e-20 * -1807217200.0 = -5.0319786e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111101001011000111100101001100;
		b = 32'b00010100001111100101010011011111;
		correct = 32'b01101000011001111111101100100010;
		#400 //0.042107865 * 9.6092865e-27 = 4.381997e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100110010000101110111000001001;
		b = 32'b10011011100101111010000010110101;
		correct = 32'b11001010001001001000110111101110;
		#400 //6.762987e-16 * -2.508471e-22 = -2696059.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011000101001110010011001101010;
		b = 32'b01110011001110010100101011101011;
		correct = 32'b10100100111001101110111100101001;
		#400 //-1470267400000000.0 * 1.4680396e+31 = -1.0015175e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000001100011010011011000000101;
		b = 32'b11101100010011001001100101000000;
		correct = 32'b00010100101100001011000000000000;
		#400 //-17.651377 * -9.893783e+26 = 1.7840878e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000100100111100000000100001110;
		b = 32'b00110010100001011110101001101000;
		correct = 32'b11010001100101110000011000111101;
		#400 //-1264.033 * 1.5589833e-08 = -81080590000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100101011000111011000010001000;
		b = 32'b01011101110110010101000001001111;
		correct = 32'b00000111000001100001110010001011;
		#400 //1.9748923e-16 * 1.9573878e+18 = 1.0089428e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110110011001111001011000011111;
		b = 32'b00001000001110001000001111111011;
		correct = 32'b01101101101000001010011101001001;
		#400 //3.4509064e-06 * 5.552563e-34 = 6.2149796e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000101101010110111100110001101;
		b = 32'b11011011111001101111110001111011;
		correct = 32'b00101001001111100000101101000011;
		#400 //-5487.194 * -1.300337e+17 = 4.2198243e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111000000001001011000110111110;
		b = 32'b11100011101111110001010000100011;
		correct = 32'b01010011101100011100011101100010;
		#400 //-1.0765441e+34 * -7.049558e+21 = 1527108600000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111011001110100001001110010100;
		b = 32'b10001110000000001111010001110110;
		correct = 32'b01101100101110001011001011010101;
		#400 //-0.0028393017 * -1.5894922e-30 = 1.7862949e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110000010111000001100011010010;
		b = 32'b00110111110101000100111001101111;
		correct = 32'b11111000000001001011001001101100;
		#400 //-2.7246683e+29 * 2.5308893e-05 = -1.0765656e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000010111010000100111101100100;
		b = 32'b01110110100100111000100101101000;
		correct = 32'b00001011110010011000110000111000;
		#400 //116.15506 * 1.4962003e+33 = 7.763336e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111001110110000001010001001100;
		b = 32'b10111101010011010010001110101001;
		correct = 32'b10111100000001101101001110000001;
		#400 //0.00041213853 * -0.050082836 = -0.008229137
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100101111110100011111001001100;
		b = 32'b01100110000010111000100010001001;
		correct = 32'b00111111011001011000111100100001;
		#400 //1.477176e+23 * 1.647319e+23 = 0.8967152
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111000011010111011100000001101;
		b = 32'b01110110110101100101000101100110;
		correct = 32'b11000001000011001100100000010111;
		#400 //-1.9123793e+34 * 2.1734424e+33 = -8.79885
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010000110110010011000000111101;
		b = 32'b01010111111100111010001000000010;
		correct = 32'b00111000011001000011011010010110;
		#400 //29150538000.0 * 535754300000000.0 = 5.4410273e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111011010101111110011010001111;
		b = 32'b11110001111111100011011100000101;
		correct = 32'b01001000110110010110101010101010;
		#400 //-1.1210201e+36 * -2.5176226e+30 = 445269.3
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011001111000110100111111000000;
		b = 32'b10110110011000000011100000110010;
		correct = 32'b11100011000000011100001111100000;
		#400 //7997813000000000.0 * -3.341131e-06 = -2.3937443e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111100101101000101011100010111;
		b = 32'b11100101011000001000111100111100;
		correct = 32'b01010110110011011001011011101101;
		#400 //-7.4910386e+36 * -6.627827e+22 = 113024050000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011000010100001110010111100101;
		b = 32'b00010001111001111101010100110101;
		correct = 32'b01000101111001101010110010100100;
		#400 //2.6999437e-24 * 3.6576773e-28 = 7381.58
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011111010011101011000011110001;
		b = 32'b01100011110111010011001101100110;
		correct = 32'b00111010111011110011010100110000;
		#400 //1.4893669e+19 * 8.160868e+21 = 0.0018250104
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101011010110110110011011010111;
		b = 32'b10111111010001010111101000000111;
		correct = 32'b00101011100011100011011000011010;
		#400 //-7.794715e-13 * -0.77139324 = 1.0104723e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101111000011000111010111010100;
		b = 32'b01101000001011001101100110000101;
		correct = 32'b00000110010100000000011110001011;
		#400 //1.2774787e-10 * 3.2650382e+24 = 3.9125994e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010001011101101100001101000000;
		b = 32'b00011111010001100110110001100100;
		correct = 32'b10110001100111110010111011010111;
		#400 //-1.9466144e-28 * 4.201779e-20 = -4.632834e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111011111000001100101100010001;
		b = 32'b01110101101000111110001001010110;
		correct = 32'b00000101101011111001001010001010;
		#400 //0.006860145 * 4.154956e+32 = 1.6510751e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100110111000111110010000110101;
		b = 32'b01100010001000000110011010010010;
		correct = 32'b00000100001101011101101110010101;
		#400 //1.5813145e-15 * 7.397175e+20 = 2.1377275e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010001111111001110110010010110;
		b = 32'b00101101010101011000110000010101;
		correct = 32'b01100100000101111001101000111111;
		#400 //135787630000.0 * 1.2138753e-11 = 1.1186292e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010000101010010110100110000101;
		b = 32'b01010101001000111010111001001111;
		correct = 32'b00111011000001000111101101011111;
		#400 //22738119000.0 * 11248065000000.0 = 0.0020215136
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010111111000111001101110010101;
		b = 32'b11101110111010110101011110000000;
		correct = 32'b00101000011101111001011001001001;
		#400 //-500514720000000.0 * -3.641738e+28 = 1.3743842e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011000011100111110000010100110;
		b = 32'b01110111101111100110111100000110;
		correct = 32'b00100000001000111110110000011011;
		#400 //1072584700000000.0 * 7.724908e+33 = 1.3884758e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001111111100110011110110001011;
		b = 32'b01111001101010010110110111110010;
		correct = 32'b00010101101101111100001100101110;
		#400 //8161793500.0 * 1.0996602e+35 = 7.422105e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101100001010101011110000011011;
		b = 32'b01000111110000110111011110011100;
		correct = 32'b00100011110111111001101110111101;
		#400 //2.4262873e-12 * 100079.22 = 2.4243666e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011100011100011011100000010000;
		b = 32'b00110001101000010010111000011000;
		correct = 32'b11101010001111111111010110011101;
		#400 //-2.721514e+17 * 4.690957e-09 = -5.8016177e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010000011110000100110001101111;
		b = 32'b00111011100011001111110101101100;
		correct = 32'b01010100011000010110110000000001;
		#400 //16663035000.0 * 0.004302671 = 3872718600000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000110100111100011101001000110;
		b = 32'b10111000110010111001111010010111;
		correct = 32'b11001101010001101110111001100100;
		#400 //20253.137 * -9.709334e-05 = -208594500.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011110111000111011010100101000;
		b = 32'b10011001000101101100010111010011;
		correct = 32'b11000101010000010101000010001011;
		#400 //2.4109484e-20 * -7.7947685e-24 = -3093.034
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000110110010100001011100000;
		b = 32'b00010100000101100011111110100111;
		correct = 32'b11011100001110010001011011100110;
		#400 //-1.5807835e-09 * 7.585618e-27 = -2.0839219e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100101000000000000011100100000;
		b = 32'b11011100000011001101111001101011;
		correct = 32'b11001000011010001010101000000110;
		#400 //3.7787146e+22 * -1.586042e+17 = -238248.1
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100010100111110011010111010001;
		b = 32'b11101011101101111111001011100101;
		correct = 32'b10110110010111011001001001001111;
		#400 //1.4684551e+21 * -4.4476092e+26 = -3.301673e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110100111000010010110101101011;
		b = 32'b01100101100011000011111000101101;
		correct = 32'b01001110110011011000010100011100;
		#400 //1.4272314e+32 * 8.278478e+22 = 1724026400.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110101000001010100000100001100;
		b = 32'b00011101111110111101010010110000;
		correct = 32'b11010110100001110111010111001110;
		#400 //-4.9641017e-07 * 6.665906e-21 = -74470020000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101010110100011000101111000010;
		b = 32'b00011100111111110110100011001110;
		correct = 32'b11001101010100100000011111001110;
		#400 //-3.7222834e-13 * 1.6901576e-21 = -220232930.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101110110101100111101001110001;
		b = 32'b11011100001101001001011010111101;
		correct = 32'b01010010000110000000010101000110;
		#400 //-3.3188907e+28 * -2.0332494e+17 = 163230880000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101110100000010101010011100110;
		b = 32'b01000100001000001100001001011110;
		correct = 32'b00101001110011011111010000001100;
		#400 //5.881322e-11 * 643.037 = 9.146164e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011110101111111110000000110111;
		b = 32'b01111010000110001011010100001111;
		correct = 32'b10100100001000001101010011010000;
		#400 //-6.9130557e+18 * 1.9822536e+35 = -3.487473e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011010000000100011100110001010;
		b = 32'b11001011011111110011100111011011;
		correct = 32'b11001110000000101001111010100100;
		#400 //9163753000000000.0 * -16726491.0 = -547858700.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011011000010101001111011010100;
		b = 32'b01000011110110001110101100011100;
		correct = 32'b10010110101000111001100001100101;
		#400 //-1.1466413e-22 * 433.8368 = -2.6430245e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001010000001110111011100000111;
		b = 32'b10001000000000001111011110011010;
		correct = 32'b01000001100001100111001011110011;
		#400 //-6.5224e-33 * -3.8809653e-34 = 16.806128
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110111011101010011100111000110;
		b = 32'b01100101000010101101101001101011;
		correct = 32'b00010001111000100000111011011110;
		#400 //1.4616589e-05 * 4.098223e+22 = 3.5665676e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111101111111111011011110100100;
		b = 32'b11100010110001111100000111111100;
		correct = 32'b11011010101000111101101110001010;
		#400 //4.2488332e+37 * -1.84244e+21 = -2.3060903e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011110111000111100101100010010;
		b = 32'b00000101001010000101000111011111;
		correct = 32'b11011001001011010011101000011101;
		#400 //-2.4118548e-20 * 7.9143594e-36 = -3047441700000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011010100100111101100111001101;
		b = 32'b10000101000110010111010011001000;
		correct = 32'b11010100111101101010011000100000;
		#400 //6.114965e-23 * -7.215475e-36 = -8474792600000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111010011101011110111010100000;
		b = 32'b01101011111111001101001000111111;
		correct = 32'b01001101111110010000011000110100;
		#400 //3.1923816e+35 * 6.1128433e+26 = 522241660.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100101010000101111110000001010;
		b = 32'b01011010010101000000110101010000;
		correct = 32'b00001010011010110110010100110001;
		#400 //1.6912212e-16 * 1.4921833e+16 = 1.13338704e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110101010000101101110101011111;
		b = 32'b11111101001110110100000011110110;
		correct = 32'b00110111100001010011001111011101;
		#400 //-2.470204e+32 * -1.5556433e+37 = 1.5878986e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000000001010100011110110100100;
		b = 32'b11011010101110101101001011110110;
		correct = 32'b00100100111010010100011011000000;
		#400 //-2.6600122 * -2.629315e+16 = 1.011675e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101100100011111011101001000100;
		b = 32'b10101001010100001011110111000111;
		correct = 32'b11000010101100000100010001101101;
		#400 //4.084984e-12 * -4.6349883e-14 = -88.133644
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101111001100100100111011100101;
		b = 32'b01001110001000110001001010001101;
		correct = 32'b00100000100010111111010101111100;
		#400 //1.6217035e-10 * 683975500.0 = 2.3709964e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111011111011010011101000000100;
		b = 32'b11001001001000100001001000000111;
		correct = 32'b10110010001110110101101101011100;
		#400 //0.007239582 * -663840.44 = -1.0905605e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111001010101001011000010110011;
		b = 32'b11111110101110010011110001100101;
		correct = 32'b00111010000100101111100010100010;
		#400 //-6.9021926e+34 * -1.2311038e+38 = 0.0005606507
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001110110101011100110010111001;
		b = 32'b10000000100010010000100010111001;
		correct = 32'b11001101110001111011010001101101;
		#400 //5.2705695e-30 * -1.2584592e-38 = -418811300.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111001101010010111111011100101;
		b = 32'b11000010100111100011001010011101;
		correct = 32'b00110110100010010010010000110000;
		#400 //-0.00032328736 * -79.098854 = 4.087131e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010111101111111100001011010010;
		b = 32'b00101111110100100010010001001110;
		correct = 32'b01100111011010011001101110101001;
		#400 //421686940000000.0 * 3.8224574e-10 = 1.1031828e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110111000000000001011011111010;
		b = 32'b11110000000001100001111010011100;
		correct = 32'b10000110011101000111110110011001;
		#400 //7.634744e-06 * -1.6603198e+29 = -4.5983574e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010001001011011100000010100001;
		b = 32'b11101010000011100001101001100110;
		correct = 32'b00100110100111001000001000011111;
		#400 //-46641320000.0 * -4.2948032e+25 = 1.0859944e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111011010001000011001001011110;
		b = 32'b11001110100001000000000111010000;
		correct = 32'b11101100001111100011110110111110;
		#400 //1.01871175e+36 * -1107355600.0 = -9.199499e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111000001001000101010110111;
		b = 32'b10001100011010011111001001001100;
		correct = 32'b01101010000100010000100101000111;
		#400 //-7.90011e-06 * -1.8022581e-31 = 4.3834514e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010111010000010010011100111110;
		b = 32'b10100001010000110110000111000101;
		correct = 32'b01110101011111010001010001110111;
		#400 //-212374290000000.0 * -6.6197967e-19 = 3.2081694e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101100110100110010001010000011;
		b = 32'b10110011011111101100101001010011;
		correct = 32'b11111000110101000010001100100001;
		#400 //2.0419706e+27 * -5.9322996e-08 = -3.4421232e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011011001011110110110001101101;
		b = 32'b11101001010110100101110011101001;
		correct = 32'b10110001010011011010100011011001;
		#400 //4.9377336e+16 * -1.6499037e+25 = -2.9927405e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001111011000110100001111011011;
		b = 32'b00011000010000101111110000101101;
		correct = 32'b00110110100101010011000011001000;
		#400 //1.12050326e-29 * 2.5201229e-24 = 4.446225e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100010100000111011111111001110;
		b = 32'b11010001000111000110101101001100;
		correct = 32'b11010000110101111001111111100011;
		#400 //1.2151722e+21 * -41988440000.0 = -28940638000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011111001110011101101000100001;
		b = 32'b01001000011111111110011101001010;
		correct = 32'b01010110001110011110110000010011;
		#400 //1.3392053e+19 * 262045.16 = 51105896000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000001101010001101011100110101;
		b = 32'b11100010000100101001001101001010;
		correct = 32'b10011111000100110111000110010011;
		#400 //21.105082 * -6.759595e+20 = -3.1222407e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111111011111011111010011010111;
		b = 32'b00000111101000110100111100110111;
		correct = 32'b01110111010001110000110001001011;
		#400 //0.9920172 * 2.4572072e-34 = 4.0371735e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010010100101100100011100010;
		b = 32'b00110001110011011101011111001001;
		correct = 32'b11001000000000110001001010101110;
		#400 //-0.0008040798 * 5.990817e-09 = -134218.72
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001000001110101010100011110000;
		b = 32'b01101010011010001111101111110111;
		correct = 32'b10011101010011010001100101110101;
		#400 //-191139.75 * 7.0415165e+25 = -2.7144685e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100100101111011010010011101001;
		b = 32'b01100001101001000011100001110100;
		correct = 32'b01000010100100111101000011110011;
		#400 //2.7986541e+22 * 3.7866674e+20 = 73.908104
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011011111101011001001111101100;
		b = 32'b10000100010110000000100001010001;
		correct = 32'b11010111000100011000000101110110;
		#400 //4.0627442e-22 * -2.5394497e-36 = -159985220000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001100111110110010110011100101;
		b = 32'b00101001100000011100110011110010;
		correct = 32'b11100010111101111011000011101101;
		#400 //-131688230.0 * 5.764303e-14 = -2.2845473e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100010010001000111010001010110;
		b = 32'b11010100110000011100001000101111;
		correct = 32'b11001101000000011100011111101101;
		#400 //9.059862e+20 * -6657492400000.0 = -136085200.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010101111110010101110111000011;
		b = 32'b00110011111010000000000000010110;
		correct = 32'b01100001100010011001010011001000;
		#400 //34272637000000.0 * 1.08033575e-07 = 3.172406e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011010000110010111001110011100;
		b = 32'b00100100110001111110010010110110;
		correct = 32'b10110100110001001000010111010110;
		#400 //-3.1733047e-23 * 8.6689944e-17 = -3.6605223e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011001111111001010101011110010;
		b = 32'b10100011001000111010101010110000;
		correct = 32'b00110110010001011001101100001011;
		#400 //-2.6125234e-23 * -8.872392e-18 = 2.9445534e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110011100100100111001001101101;
		b = 32'b10011011110111001111000000111011;
		correct = 32'b01010111001010011010111111101110;
		#400 //-6.819469e-08 * -3.6551192e-22 = 186573080000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000010111011101001100101000001;
		b = 32'b00111101010000010101011000111011;
		correct = 32'b11000101000111011111011101000101;
		#400 //-119.299324 * 0.047201376 = -2527.4543
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011110011111000011101100011101;
		b = 32'b11010011100010100100000000101111;
		correct = 32'b11001010011010011000011101101111;
		#400 //4.5437882e+18 * -1187564600000.0 = -3826139.8
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000110001010111010111101010110;
		b = 32'b10110000011110011010011001011111;
		correct = 32'b00010101001100000000110101001001;
		#400 //-3.2290342e-35 * -9.08221e-10 = 3.5553397e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100111000111001110010001110111;
		b = 32'b01001000011010000010101110111110;
		correct = 32'b10011110001011001111111011001011;
		#400 //-2.17732e-15 * 237742.97 = -9.158294e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111100100111110000010010010;
		b = 32'b10110000000111010000110000110100;
		correct = 32'b11010110111100010000110100101101;
		#400 //75713.14 * -5.713361e-10 = -132519450000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011111100110111101001111100000;
		b = 32'b00101110011000010001010011010100;
		correct = 32'b00110000101100010011101110101111;
		#400 //6.599557e-20 * 5.1177576e-11 = 1.2895408e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011100111001100101100100100001;
		b = 32'b01110010101110110010011101001110;
		correct = 32'b10101001100111011000101011001000;
		#400 //-5.1869794e+17 * 7.413915e+30 = -6.996275e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011000000110100100111101111111;
		b = 32'b10110000110011011001111010101010;
		correct = 32'b01100110110000000001111010000000;
		#400 //-678664900000000.0 * -1.4960808e-09 = 4.536285e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000111111101100010100011110000;
		b = 32'b10000011100001011000100010000000;
		correct = 32'b11000011111010111111010110110110;
		#400 //3.7038027e-34 * -7.848376e-37 = -471.91962
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100011000000101011101001000101;
		b = 32'b01100000111101010011111001011010;
		correct = 32'b01000001100010000111011000011100;
		#400 //2.411499e+21 * 1.4137329e+20 = 17.05767
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011001000010001010101001111100;
		b = 32'b01001101001001000100101110011110;
		correct = 32'b00001011010101001111001011011101;
		#400 //7.065464e-24 * 172276200.0 = 4.1012425e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010100100101111011101100111001;
		b = 32'b00111110011100010000010011010110;
		correct = 32'b01010101101000010010100110011110;
		#400 //5213449000000.0 * 0.23537001 = 22150015000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101000001011011111111000010000;
		b = 32'b01011000110111110100100101000011;
		correct = 32'b01001110110001110111101111110100;
		#400 //3.286624e+24 * 1964046000000000.0 = 1673394700.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110000110101001100111111100101;
		b = 32'b01100100101000010001010101010010;
		correct = 32'b11001011101010010001101011010001;
		#400 //-5.268972e+29 * 2.3771697e+22 = -22164898.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110100111101011111100111111000;
		b = 32'b11001111001100011001011100000100;
		correct = 32'b11100101001100010100101001010111;
		#400 //1.5590609e+32 * -2979464200.0 = -5.2326887e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111110110010111110111101010010;
		b = 32'b11101001111010111001000100110110;
		correct = 32'b11010100010111011001111110110110;
		#400 //1.3553795e+38 * -3.5597913e+25 = -3807469000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101001101001011001011001101101;
		b = 32'b10011010000110111001011010011100;
		correct = 32'b11001111000010000011100111101011;
		#400 //7.353567e-14 * -3.217491e-23 = -2285497000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000001001100110001001011000111;
		b = 32'b11101010111000101100111010000011;
		correct = 32'b10010101110010100001111101101001;
		#400 //11.192084 * -1.3709623e+26 = -8.1636707e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000010000001100100001001010100;
		b = 32'b11011101100011011100111001001011;
		correct = 32'b10100011111100100110000001000001;
		#400 //33.564774 * -1.2772734e+18 = -2.6278458e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011000110110110101100111000011;
		b = 32'b01111111111000000111001111111001;
		correct = 32'b01111111111000000111001111111001;
		#400 //-1929428600000000.0 * nan = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101011001101110000011011011100;
		b = 32'b10110011110111010001010111011111;
		correct = 32'b10110110110100111110111001010111;
		#400 //6.502418e-13 * -1.0295093e-07 = -6.3160364e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001110001000111010110001111010;
		b = 32'b01110011101001001010111000111111;
		correct = 32'b00011001111111100110111101001011;
		#400 //686497400.0 * 2.609469e+31 = 2.6307935e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110001011111010010011010100111;
		b = 32'b10111111000100010011010110000111;
		correct = 32'b10110001110111110010011001000001;
		#400 //3.6838317e-09 * -0.567223 = -6.494503e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111011001001101011100101101010;
		b = 32'b00100010100111110001000000001010;
		correct = 32'b01011000000001100010101001011001;
		#400 //0.0025440105 * 4.311402e-18 = 590065760000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001100011100011011010110110011;
		b = 32'b00001010000010100100001100111010;
		correct = 32'b11000001110111111100010011001101;
		#400 //-1.8620643e-31 * 6.657102e-33 = -27.971094
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111101000000111000001100010110;
		b = 32'b00100101101111011100100110001010;
		correct = 32'b11010110101100010110010011010001;
		#400 //-0.032107435 * 3.2922842e-16 = -97523280000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010010010100101101110101111100;
		b = 32'b00111101111011101001101100011000;
		correct = 32'b01010011111000100011110010110000;
		#400 //226414760000.0 * 0.116506755 = 1943361600000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110001000101110011111101100111;
		b = 32'b11000100010110001001110000100111;
		correct = 32'b11101100001100101100000001110000;
		#400 //7.489422e+29 * -866.4399 = -8.643902e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011101110100011000001100011000;
		b = 32'b10101101101011001011110001101111;
		correct = 32'b11101111100110110100000001100111;
		#400 //1.8871171e+18 * -1.9637817e-11 = -9.609607e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111110101010000000110101011000;
		b = 32'b01111010000001111110001101110100;
		correct = 32'b01000100000111100100101111100111;
		#400 //1.1168979e+38 * 1.7639334e+35 = 633.186
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101001101011010101110000000011;
		b = 32'b01001001100001101010001001101100;
		correct = 32'b01011111101001001101000100010010;
		#400 //2.6197335e+25 * 1102925.5 = 2.3752587e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000010101110001111101101101010;
		b = 32'b11001001110100110001111110000011;
		correct = 32'b00111000011000000100110101101001;
		#400 //-92.49104 * -1729520.4 = 5.3477856e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110111011001011101010110110010;
		b = 32'b11101111110001111101101101000111;
		correct = 32'b01000111000100110011001100100111;
		#400 //-4.6616025e+33 * -1.2370521e+29 = 37683.152
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100100000000010101010101110011;
		b = 32'b01010110111001101100110111011001;
		correct = 32'b00001100100011110111001111011110;
		#400 //2.8044794e-17 * 126885890000000.0 = 2.2102374e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110100110001000000111010101111;
		b = 32'b01010000000101000111010001101000;
		correct = 32'b00100100001010010000101100110011;
		#400 //3.651853e-07 * 9962627000.0 = 3.665552e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100111011011111111110110011011;
		b = 32'b10111101010100000110000100000101;
		correct = 32'b10101001100100110110101011111111;
		#400 //3.3305393e-15 * -0.050873775 = -6.546672e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010111000110100010101001010001;
		b = 32'b11110110001101110010110110110101;
		correct = 32'b10100000010101110111001111100110;
		#400 //169506540000000.0 * -9.2882556e+32 = -1.8249556e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000011101100000101000110010000;
		b = 32'b10000101101000001010111101011011;
		correct = 32'b01111101100011000111010000011110;
		#400 //-352.6372 * -1.5110743e-35 = 2.3336854e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101100000010100100100000010000;
		b = 32'b01101000110000111000001001010101;
		correct = 32'b11000010101101010001000011101001;
		#400 //-6.686883e+26 * 7.3861253e+24 = -90.53303
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000001011000001011011101001110;
		b = 32'b10111100100011010011011001000010;
		correct = 32'b01000100010010111011000011111101;
		#400 //-14.044752 * -0.017237786 = 814.76544
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110000001001000000101000100011;
		b = 32'b00010101101110011000100101010000;
		correct = 32'b01011001111000100101011011001111;
		#400 //5.967726e-10 * 7.4937546e-26 = 7963599000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011000011111010101011111011111;
		b = 32'b00010010000011100011010111001110;
		correct = 32'b01000101111001000000011100111011;
		#400 //3.2743847e-24 * 4.487362e-28 = 7296.904
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000000010110111011111011101000;
		b = 32'b10001101110100111001010000001001;
		correct = 32'b11110010000001001111000011101110;
		#400 //3.433527 * -1.3039517e-30 = -2.6331704e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010001111010110001111011110011;
		b = 32'b10100100100110111101001001000100;
		correct = 32'b01101100110000010010010000010010;
		#400 //-126229570000.0 * -6.757674e-17 = 1.8679442e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001001111101010111000100100100;
		b = 32'b01000010001101000001011101111111;
		correct = 32'b00000111001011100111001010010011;
		#400 //5.9088e-33 * 45.022945 = 1.3123975e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111001011100011110001001000111;
		b = 32'b11000001110011100011110011000010;
		correct = 32'b00110111000101100001111110110011;
		#400 //-0.00023067846 * -25.779667 = 8.948077e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011001100100100110000110011110;
		b = 32'b00001001111111010010000000011001;
		correct = 32'b11001111000101000000101100110000;
		#400 //-1.5135473e-23 * 6.093772e-33 = -2483761200.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001000100111001101111110110111;
		b = 32'b11000111111001110000110001101111;
		correct = 32'b11000000001011011101000010100110;
		#400 //321277.72 * -118296.87 = -2.71586
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101100011011100101100001000001;
		b = 32'b01110010111110111111001101010100;
		correct = 32'b10111000111100100010110011110010;
		#400 //-1.15256445e+27 * 9.9807876e+30 = -0.00011547831
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011011111101100100101011100010;
		b = 32'b00010110011111111111111101001001;
		correct = 32'b01000100111101100100101110010010;
		#400 //4.0745678e-22 * 2.067929e-25 = 1970.3616
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100110101100110001100101100000;
		b = 32'b10010100101010000111101111010100;
		correct = 32'b11010001100010000001000010010001;
		#400 //1.2427498e-15 * -1.7012506e-26 = -73049190000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000010111000011001101000111100;
		b = 32'b11100010101001100111001010011101;
		correct = 32'b00011111101011010111110110011010;
		#400 //-112.80124 * -1.5352091e+21 = 7.347614e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110011010000000101101000110111;
		b = 32'b10101101011110000000001011101001;
		correct = 32'b01000101010001101000110001011000;
		#400 //-4.4785534e-08 * -1.4097814e-11 = 3176.7715
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001110001011100100111011001001;
		b = 32'b11101100000011010101111100001000;
		correct = 32'b10100001100111011101001001000010;
		#400 //731099700.0 * -6.8362925e+26 = -1.0694389e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011001101011110110111011101001;
		b = 32'b10100100001100111100101010000011;
		correct = 32'b10110100111110011100101110000110;
		#400 //1.8139372e-23 * -3.8985972e-17 = -4.6527947e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001011111010101110100000001101;
		b = 32'b00000010011110101101000010111111;
		correct = 32'b01001000111011111100001100011110;
		#400 //9.048267e-32 * 1.8427006e-37 = 491032.94
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100000110110111000001001010000;
		b = 32'b10011010100010111101011101011111;
		correct = 32'b01000101110010001110101111110111;
		#400 //-3.7186277e-19 * -5.7837003e-23 = 6429.4956
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101010000011101000010111011101;
		b = 32'b01000100001110001101111010101100;
		correct = 32'b00100101010001010101110000011010;
		#400 //1.2658577e-13 * 739.47925 = 1.7118231e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001101011011110011000011110000;
		b = 32'b11000111010101001001111111011101;
		correct = 32'b10000101100011111111111001000000;
		#400 //7.3706467e-31 * -54431.863 = -1.3541052e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100101100011100011101100111001;
		b = 32'b01100001011010001110110111101101;
		correct = 32'b00000011100111000101000110010111;
		#400 //2.4673204e-16 * 2.6854931e+20 = 9.187588e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001100101001011010110101010010;
		b = 32'b00101110011011000110011111010000;
		correct = 32'b10011101101100110110100011000000;
		#400 //-2.5526589e-31 * 5.375239e-11 = -4.7489214e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011010000000000001101101001100;
		b = 32'b11110111000110011101000001011001;
		correct = 32'b00100010010101010011011011010101;
		#400 //-9014703000000000.0 * -3.1197157e+33 = 2.889591e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100100011100001101100100001111;
		b = 32'b10011110001101111010001011100001;
		correct = 32'b01000101101001111110000011010100;
		#400 //-5.222556e-17 * -9.721622e-21 = 5372.1035
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100100010001110111111110100001;
		b = 32'b10010011110010011100100101011101;
		correct = 32'b01001111111111010001100011100110;
		#400 //-4.3259352e-17 * -5.0938093e-27 = 8492535000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001010110011001101100110101010;
		b = 32'b11001110100101111011101010000111;
		correct = 32'b10111011101011001101000001100011;
		#400 //6712533.0 * -1272791900.0 = -0.005273865
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010110101010010010011101010001;
		b = 32'b10111111000100010100111001101001;
		correct = 32'b10010111000101010000000111001101;
		#400 //2.7328235e-25 * -0.5676027 = -4.814677e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111101101100011000101110010001;
		b = 32'b01110101011001001100010101110100;
		correct = 32'b10000111110001101010110101000111;
		#400 //-0.08669198 * 2.9000208e+32 = -2.9893572e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011001011011011011011101001011;
		b = 32'b00110001010110001110111100100011;
		correct = 32'b11100111100011000100001100011100;
		#400 //-4181944000000000.0 * 3.156807e-09 = -1.3247385e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010101010001101110010011100000;
		b = 32'b00111011010110000011110110100110;
		correct = 32'b00011001011010110111011010111001;
		#400 //4.0166332e-26 * 0.003299573 = 1.2173191e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000010110110000011010100000011;
		b = 32'b10110110001110101010001100100000;
		correct = 32'b00001100000101000100011110011001;
		#400 //-3.1768775e-37 * -2.781111e-06 = 1.1423051e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101010111000000000100100101001;
		b = 32'b01100111111110101101001011000010;
		correct = 32'b10000010011001001010100011011110;
		#400 //-3.979675e-13 * 2.3689588e+24 = -1.6799257e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100101111010000000111010000110;
		b = 32'b11111110110010000110001011110000;
		correct = 32'b00100110100101000011101011011001;
		#400 //-1.3698212e+23 * -1.3317966e+38 = 1.0285514e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110001011001001110000111000010;
		b = 32'b11110010010111001011001011101100;
		correct = 32'b00111110100001001011111011110100;
		#400 //-1.1333681e+30 * -4.3713923e+30 = 0.25926936
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001011111010101011111110001101;
		b = 32'b00100110010001000101001000010110;
		correct = 32'b10100101000110010000110111111001;
		#400 //-9.0421735e-32 * 6.811241e-16 = -1.3275369e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010011011010100010101011000110;
		b = 32'b01111010101110101011111100000110;
		correct = 32'b10011000001000001000000011011011;
		#400 //-1005739970000.0 * 4.848208e+35 = -2.074457e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001111101011010101000101011100;
		b = 32'b00101001000010111010001011111000;
		correct = 32'b00100110000111101101111111011000;
		#400 //1.7090456e-29 * 3.1005553e-14 = 5.5120627e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000111000111010011101000110101;
		b = 32'b10000001011010011100110000111000;
		correct = 32'b01000101001011000010100010000011;
		#400 //-1.1828473e-34 * -4.294186e-38 = 2754.532
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000111000000111111111010010;
		b = 32'b11001000100111100110001001110111;
		correct = 32'b00100111101101010110111001100010;
		#400 //-1.6334474e-09 * -324371.72 = 5.035727e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001010010110111011110001001110;
		b = 32'b10011000010000111101010110011110;
		correct = 32'b01110001100011111001111101000001;
		#400 //-3600147.5 * -2.5311008e-24 = 1.4223642e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100111000110011100011010010110;
		b = 32'b01001111010101100000110001110010;
		correct = 32'b10010111001101111110101000001011;
		#400 //-2.134067e-15 * 3591139800.0 = -5.9425893e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100000001101000110110101110111;
		b = 32'b11011101111010101000001100101110;
		correct = 32'b01000001110001001111010110100110;
		#400 //-5.2004714e+19 * -2.1123001e+18 = 24.619946
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110001101010100000011000110101;
		b = 32'b10110111111111110001010101000110;
		correct = 32'b11111001001010101010001010101010;
		#400 //1.6838386e+30 * -3.0408275e-05 = -5.5374355e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100000010110111001101010111010;
		b = 32'b01000010010011100010001110110000;
		correct = 32'b00011101100010000101110001100111;
		#400 //1.8601216e-19 * 51.53485 = 3.6094442e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111000010011111010000001010010;
		b = 32'b11000110101100000000111101011001;
		correct = 32'b10110001000101101111001100010010;
		#400 //4.9501956e-05 * -22535.674 = -2.1966042e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111001100011110101000001000111;
		b = 32'b10001100000000110000101101100001;
		correct = 32'b01101101000010111111101111101110;
		#400 //-0.00027334897 * -1.0095297e-31 = 2.7076863e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010011100101010101001110101001;
		b = 32'b01111010101011000010101001011110;
		correct = 32'b10011000010111100000101001001010;
		#400 //-1282707400000.0 * 4.469672e+35 = -2.8698022e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101100110001010100100001000111;
		b = 32'b01011101000001100010101100001110;
		correct = 32'b10001111001111000011011001101011;
		#400 //-5.607101e-12 * 6.042398e+17 = -9.279596e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110010000010111000000111111110;
		b = 32'b10100000100111101100110001010101;
		correct = 32'b11010000111000001110011011011011;
		#400 //8.120422e-09 * -2.6901457e-19 = -30185806000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011100111001100001110110000001;
		b = 32'b10111011111101011101010010000001;
		correct = 32'b11100000011011111010001010010010;
		#400 //5.1817348e+17 * -0.007502139 = -6.9070098e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011101011001110011010100010100;
		b = 32'b01010011010001000101100100100110;
		correct = 32'b00001001100101101011100110001001;
		#400 //3.0600036e-21 * 843309250000.0 = 3.6285663e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001001101110110001000111010000;
		b = 32'b11111010110110111010011011010100;
		correct = 32'b00001110010110100000011010110011;
		#400 //-1532474.0 * -5.7024834e+35 = 2.68738e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010111000001101100111111010100;
		b = 32'b11111011000011000100111010100100;
		correct = 32'b10011011011101011111100100101101;
		#400 //148227170000000.0 * -7.285166e+35 = -2.0346438e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000101011100001100001001011111;
		b = 32'b10110010001110000001101100111000;
		correct = 32'b01010010101001110110001101010011;
		#400 //-3852.1482 * -1.0716398e-08 = 359462960000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110110111001011000011110111;
		b = 32'b00111000111101100001111000111110;
		correct = 32'b10111101011001011000110101011111;
		#400 //-6.5771123e-06 * 0.00011735827 = -0.056043025
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011000010100101101000100110111;
		b = 32'b01111101001111000100011101110110;
		correct = 32'b10011010100011110101001010000101;
		#400 //-927184050000000.0 * 1.5641619e+37 = -5.927673e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100011101110100010100110001001;
		b = 32'b01010001001100001111110000110011;
		correct = 32'b10010010000001101010001100011001;
		#400 //-2.0183751e-17 * 47509090000.0 = -4.248398e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110101001010011101001000101011;
		b = 32'b11101010011000011001011101011111;
		correct = 32'b10001010010000001011011001001011;
		#400 //6.326324e-07 * -6.8180785e+25 = -9.278749e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010011110011111101110111110110;
		b = 32'b10001110101010101000001110001011;
		correct = 32'b11000100100111000000101000111110;
		#400 //5.2473017e-27 * -4.2034907e-30 = -1248.3201
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101101100101011101100000101000;
		b = 32'b10111011111011101000000001110010;
		correct = 32'b11110001001000001101011010001011;
		#400 //5.796823e+27 * -0.0072784955 = -7.964315e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100111110010101010000101011011;
		b = 32'b10001111111111000111100011010110;
		correct = 32'b11010111010011010111011000111001;
		#400 //5.6241205e-15 * -2.4895663e-29 = -225907650000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111000001010100011110011110101;
		b = 32'b00101101011100001010010110000101;
		correct = 32'b11001010001101010001100101110101;
		#400 //-4.058793e-05 * 1.3679173e-11 = -2967133.2
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010011000100010101001000101001;
		b = 32'b00111000010100111010010110000010;
		correct = 32'b00011010001011111100011001100101;
		#400 //1.8342081e-27 * 5.046046e-05 = 3.6349414e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001100101110111111101010001100;
		b = 32'b11010001110000010110111010011001;
		correct = 32'b00111010011110001100100001100001;
		#400 //-98554980.0 * -103848030000.0 = 0.0009490308
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001000100011000111100000111100;
		b = 32'b10111111110101011011001001111010;
		correct = 32'b11001000001010000100011011001111;
		#400 //287681.88 * -1.6695092 = -172315.23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110010110101000000011010101001;
		b = 32'b10010010000001100011011100110000;
		correct = 32'b11100000010010100011010011111110;
		#400 //2.4683077e-08 * -4.235097e-28 = -5.82822e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110000000010111111001000011110;
		b = 32'b10001100010101011100100001001100;
		correct = 32'b11100011001001111001010100001000;
		#400 //5.0911975e-10 * -1.6469198e-31 = -3.091345e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111101001010111000001010011;
		b = 32'b10110010011101110010101001100101;
		correct = 32'b11010100101010110101101000011110;
		#400 //84704.65 * -1.4386932e-08 = -5887610600000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111100001101100110011000110100;
		b = 32'b01011000111001001001001110001100;
		correct = 32'b01100010110011000100100001100001;
		#400 //3.7882838e+36 * 2010578900000000.0 = 1.8841756e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010101001000100000000100011011;
		b = 32'b01011111000101110001111100101100;
		correct = 32'b00110101100010010011011110101111;
		#400 //11132852000000.0 * 1.0889471e+19 = 1.0223501e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010001010011111000011010000011;
		b = 32'b01111101000001000100010001010011;
		correct = 32'b00010011110010001101010010101010;
		#400 //55707185000.0 * 1.0988303e+37 = 5.06968e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000101010111010010001100001011;
		b = 32'b00110101110111110111000010101101;
		correct = 32'b01001110111111010101110001110010;
		#400 //3538.1902 * 1.6647588e-06 = 2125347100.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000000110101110000011010100;
		b = 32'b00100011111000110110111101111000;
		correct = 32'b11001011101011100101010001111110;
		#400 //-5.6344374e-10 * 2.4658598e-17 = -22849788.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000110000101111111010010110111;
		b = 32'b00101000101110100010110100011011;
		correct = 32'b01011100110100001111001000011001;
		#400 //9725.179 * 2.066971e-14 = 4.7050387e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100000011001100001101010011101;
		b = 32'b11010110010001111110111001011001;
		correct = 32'b11001001100100110101000100111100;
		#400 //6.632295e+19 * -54956627000000.0 = -1206823.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001001111111000110010100000000;
		b = 32'b00101100111110000110100001100111;
		correct = 32'b01011100100000100000110111100101;
		#400 //2067616.0 * 7.060175e-12 = 2.928562e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110111010101010110110101000100;
		b = 32'b01000000100100010001101100010010;
		correct = 32'b00110110001111000100010001011111;
		#400 //1.272123e-05 * 4.5345545 = 2.805398e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001000101001000011110011010100;
		b = 32'b01001000100011110000101011000001;
		correct = 32'b10111111100100101111011101111011;
		#400 //-336358.62 * 292950.03 = -1.1481775
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011111000001110110010101011110;
		b = 32'b11011101010110110011000001111101;
		correct = 32'b00000001000111100010001001100011;
		#400 //-2.867121e-20 * -9.871413e+17 = 2.9044688e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001110010001101101100111100100;
		b = 32'b00110100000111000111111001110111;
		correct = 32'b00011001101000101010010100010110;
		#400 //2.4510295e-30 * 1.457464e-07 = 1.6817085e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110110010110110100010010011010;
		b = 32'b11011100111010010110001001010101;
		correct = 32'b01011000111100001000010000010110;
		#400 //-1.1118207e+33 * -5.255343e+17 = 2115600800000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010111001011101101110100000111;
		b = 32'b01000010111101010001001000001001;
		correct = 32'b01010011101101101010100101110000;
		#400 //192264330000000.0 * 122.535225 = 1569053500000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000111111011101100111101010011;
		b = 32'b00011111011100001011011110101110;
		correct = 32'b11100111111111011111100010100100;
		#400 //-122270.65 * 5.0973913e-20 = -2.3986907e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010001010001011011111010000001;
		b = 32'b01000001011000010101111000101001;
		correct = 32'b10001111011000001001111100101000;
		#400 //-1.5599263e-28 * 14.085488 = -1.1074705e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010100011011110111000010001110;
		b = 32'b00000001110101100110111000100100;
		correct = 32'b01010010000011101110110111001100;
		#400 //1.2088614e-26 * 7.876923e-38 = 153468730000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010010111010110000011101110010;
		b = 32'b00101011001110001000101000110111;
		correct = 32'b10100111001000110000010100101001;
		#400 //-1.483242e-27 * 6.5561743e-13 = -2.2623591e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010000000101000110010011001111;
		b = 32'b00110111101011001111010010110000;
		correct = 32'b01010111110110111010010100000100;
		#400 //9958538000.0 * 2.061794e-05 = 483003570000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001010100011110101010111100101;
		b = 32'b01011111111101011011011011100100;
		correct = 32'b10101010000101010101010111100110;
		#400 //-4696818.5 * 3.541118e+19 = -1.326366e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100110111011000110110110101000;
		b = 32'b01011101001010110111001010110111;
		correct = 32'b01001001001100001000001101010111;
		#400 //5.5825065e+23 * 7.721336e+17 = 722997.44
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111000101011001110001111000101;
		b = 32'b11110100011101001111100000001110;
		correct = 32'b11000011101101001010110011001101;
		#400 //2.8052962e+34 * -7.7633763e+31 = -361.35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010011000110110110011001101111;
		b = 32'b01101110001110001010010111100111;
		correct = 32'b10100100010101110111001100110111;
		#400 //-667438500000.0 * 1.4286451e+28 = -4.6718284e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010010101101100001110101011010;
		b = 32'b00000011110001100111100011010111;
		correct = 32'b11001110011010101110011011000000;
		#400 //-1.14930505e-27 * 1.16651375e-36 = -985247740.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011100111111011001001101110;
		b = 32'b01100101111100110100000011001100;
		correct = 32'b10100101001010000001000010111110;
		#400 //-20931804.0 * 1.4359129e+23 = -1.457735e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011111100100000111100000110011;
		b = 32'b11011011001111001001101001000000;
		correct = 32'b01000011110001000001100010010010;
		#400 //-2.0820253e+19 * -5.3086895e+16 = 392.19196
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110110000011110011010100001101;
		b = 32'b11100001100111001110100001110110;
		correct = 32'b10010011111010011010010110001111;
		#400 //2.133954e-06 * -3.6180533e+20 = -5.8980722e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100010010101000000111001000111;
		b = 32'b01000100001010011111111010000110;
		correct = 32'b11011101100111111010101111000011;
		#400 //-9.779346e+20 * 679.9769 = -1.438188e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110000011111011010100000101100;
		b = 32'b11010101000110100001001001101111;
		correct = 32'b01011010110100101011101110110011;
		#400 //-3.1401206e+29 * -10587748000000.0 = 2.9658061e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110110011111000000110100001101;
		b = 32'b01110101110111011010001001110010;
		correct = 32'b11000000000100011001000011111010;
		#400 //-1.2780503e+33 * 5.6191035e+32 = -2.2744737
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000100101101101110100010101100;
		b = 32'b10011111011001010101000110010100;
		correct = 32'b10100100110011000011000010111111;
		#400 //4.300167e-36 * -4.8560116e-20 = -8.8553476e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010101001001111000100101111101;
		b = 32'b11000101000011011010101111010010;
		correct = 32'b01001111100101110101111010101110;
		#400 //-11513059000000.0 * -2266.7388 = 5079129000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111001000110101111100001110;
		b = 32'b00001011101000100110101000100100;
		correct = 32'b01111011000000001100000100000101;
		#400 //41823.055 * 6.255983e-32 = 6.685289e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001000100110100110011100100000;
		b = 32'b10111111101010110100001101100011;
		correct = 32'b10001000011001101100110000101001;
		#400 //9.292782e-34 * -1.337994 = -6.9453096e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111001101000011010110111011010;
		b = 32'b11011000000001111100010101101111;
		correct = 32'b10100001000110000110110011001011;
		#400 //0.00030837842 * -597128160000000.0 = -5.164359e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010000101011011010000010000110;
		b = 32'b11001101000111110010010100000110;
		correct = 32'b01000011000010111010010111110001;
		#400 //-23303827000.0 * -166875230.0 = 139.64821
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100100000111101001111000001011;
		b = 32'b10110100000011000000000001101000;
		correct = 32'b10101111100100010000010100011011;
		#400 //3.4394656e-17 * -1.3038664e-07 = -2.6378974e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001110100110011011110001111100;
		b = 32'b10110100010100100001110110110001;
		correct = 32'b01011001101110110100111011110010;
		#400 //-1289633300.0 * -1.9568576e-07 = 6590328000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101000101000000100000100101101;
		b = 32'b11000001110001111110111110100011;
		correct = 32'b11100110010011010011000100000011;
		#400 //6.0542473e+24 * -24.99201 = -2.422473e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001001111101110100000000101011;
		b = 32'b10110000111000100011011110011011;
		correct = 32'b00011000100010111110011010111100;
		#400 //-5.952343e-33 * -1.6459468e-09 = 3.616364e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010010000010101001001000011110;
		b = 32'b01000111000001100001010101101101;
		correct = 32'b01001010100001000100100010010011;
		#400 //148789230000.0 * 34325.426 = 4334665.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111001100111000100011011001010;
		b = 32'b11100111010110000110011111100110;
		correct = 32'b11010001101110001101111010001000;
		#400 //1.0142926e+35 * -1.02194775e+24 = -99250930000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101110000100100011111101100100;
		b = 32'b10111100001000101011011110100101;
		correct = 32'b01110001011001100001011010100111;
		#400 //-1.1315361e+28 * -0.00993148 = 1.139343e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011110110100100110101001001011;
		b = 32'b00110100010110010101001000010000;
		correct = 32'b00101001111101111101110110011001;
		#400 //2.2278577e-20 * 2.0239554e-07 = 1.10074445e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010101001001101010011011000100;
		b = 32'b00111100001110000100110100101111;
		correct = 32'b00011000011001110111101111001010;
		#400 //3.3654988e-26 * 0.011248871 = 2.9918548e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000100001000001111110111101001;
		b = 32'b00101000110010000111101000000110;
		correct = 32'b00011010110011011001010001100001;
		#400 //1.89245e-36 * 2.225738e-14 = 8.502573e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110110110010110010000111110;
		b = 32'b10100110000100010111010110100110;
		correct = 32'b11011000001111110100110001001001;
		#400 //0.4245929 * -5.0466424e-16 = -841337450000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011000100101001100000110100111;
		b = 32'b01100101100100000100100111110101;
		correct = 32'b10110010100000111111011010010101;
		#400 //-1308475600000000.0 * 8.517313e+22 = -1.536254e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010101110001010001001001000101;
		b = 32'b01001001101000000111000011111011;
		correct = 32'b11001011100111010011100100110010;
		#400 //-27085282000000.0 * 1314335.4 = -20607588.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100011110100010000011100010000;
		b = 32'b01101111010101101110100000010000;
		correct = 32'b10110011111110001111111100111000;
		#400 //-7.711757e+21 * 6.651034e+28 = -1.1594824e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000011011100101010100100000100;
		b = 32'b11010000011000011001100111001111;
		correct = 32'b10110010100010011010110111010111;
		#400 //242.66022 * -15139814000.0 = -1.6027952e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011010110100111111101111011101;
		b = 32'b01010001011000100001101110010010;
		correct = 32'b01001000111100000000001001001000;
		#400 //2.9834073e+16 * 60695323000.0 = 491538.25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001001101111110110100010000011;
		b = 32'b00100100000101011100011001111101;
		correct = 32'b11100101001000111001010001111101;
		#400 //-1568016.4 * 3.247735e-17 = -4.8280304e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100001100111011110100010000000;
		b = 32'b11100010111100000101001011100001;
		correct = 32'b10111110001010000011010101100001;
		#400 //3.6411153e+20 * -2.2165953e+21 = -0.16426612
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011010100100110111100101101000;
		b = 32'b01010000100111110111010000111110;
		correct = 32'b10001001011011001100010001000011;
		#400 //-6.099392e-23 * 21401563000.0 = -2.8499748e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011111011100001111100010100001;
		b = 32'b11010101001111110001100001100010;
		correct = 32'b11001001101000010110100001110111;
		#400 //1.7363805e+19 * -13131965000000.0 = -1322254.9
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101010110001001110110110111011;
		b = 32'b01011010010101000110101100010010;
		correct = 32'b01001111111011010101010100011000;
		#400 //1.1903606e+26 * 1.4947605e+16 = 7963554000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010110011001001111010001100010;
		b = 32'b00111011101010111001101100011101;
		correct = 32'b01011010001010101100011010110000;
		#400 //62934567000000.0 * 0.005236997 = 1.2017301e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010101100001001111100100110111;
		b = 32'b01001011011101101000000011000111;
		correct = 32'b00001001100010100001100010110110;
		#400 //5.370757e-26 * 16154823.0 = 3.324553e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101111000100110000100010010111;
		b = 32'b00110000101100101000000010100111;
		correct = 32'b00111101110100101101111001011111;
		#400 //1.3372624e-10 * 1.298777e-09 = 0.1029632
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100111101111110101001011110110;
		b = 32'b10100001001110011110110000010011;
		correct = 32'b11000110000000111011100000010000;
		#400 //5.3103096e-15 * -6.299288e-19 = -8430.016
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100011100110000011001111000001;
		b = 32'b11011110011000001100101011010111;
		correct = 32'b01000100101011010101010100001100;
		#400 //-5.615269e+21 * -4.0494989e+18 = 1386.6577
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011100101101110010001111100000;
		b = 32'b00100011000000100110011001001100;
		correct = 32'b01111001001100111100010100100000;
		#400 //4.1239493e+17 * 7.068976e-18 = 5.8338707e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101010111010001000011000101111;
		b = 32'b11010101101110010101101110010110;
		correct = 32'b01010100101000001001001000110001;
		#400 //-1.4055223e+26 * -25475376000000.0 = 5517179600000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111111101110010000101111001111;
		b = 32'b10010000110100111100010100011110;
		correct = 32'b01101110010111111011000111010011;
		#400 //-1.4456729 * -8.352853e-29 = 1.7307533e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000110101011111100101101010001;
		b = 32'b00110001101011000111110111001001;
		correct = 32'b00010100100000100111001101110001;
		#400 //6.612643e-35 * 5.020159e-09 = 1.3172179e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011010000010010010001000001000;
		b = 32'b00001001110000011000111011000001;
		correct = 32'b11001111101101010101111101011100;
		#400 //-2.8358426e-23 * 4.6597305e-33 = -6085851000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011011010101110010100111100110;
		b = 32'b00110000111010100111101111111011;
		correct = 32'b01101001111010101110100000010100;
		#400 //6.0563188e+16 * 1.7060978e-09 = 3.5498075e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100110000100010100011011111000;
		b = 32'b11000010010000010101000100110101;
		correct = 32'b00100011010000000110001000010100;
		#400 //-5.040316e-16 * -48.329304 = 1.042911e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100101111010001101110001111011;
		b = 32'b00111100000111111100101101010001;
		correct = 32'b00101001001110101000011101100111;
		#400 //4.0394988e-16 * 0.009753064 = 4.141774e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000110000110101011100000011010;
		b = 32'b11000110111111100101000010001111;
		correct = 32'b10111110100110111011111010010101;
		#400 //9902.025 * -32552.28 = -0.3041884
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011011001011001000011000111111;
		b = 32'b00101110011100000011010110011001;
		correct = 32'b10101100001101111101110110011010;
		#400 //-1.4270884e-22 * 5.4617286e-11 = -2.6128878e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100010001111110110011100000100;
		b = 32'b11010100010101101100101000011110;
		correct = 32'b10001101011001000010000000110000;
		#400 //2.5939863e-18 * -3690055900000.0 = -7.029667e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011001111100000110010000010111;
		b = 32'b00100101101011001101111010111011;
		correct = 32'b11110011101100011111111011001000;
		#400 //-8458005500000000.0 * 2.9988172e-16 = -2.8204471e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001111001101110110100001101001;
		b = 32'b00001001011001011110011000100001;
		correct = 32'b01000101010011000011101100001100;
		#400 //9.042705e-30 * 2.7673078e-33 = 3267.6904
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101101110010000111101000011010;
		b = 32'b00011000111110001010000011001011;
		correct = 32'b01010100010011100110101111010001;
		#400 //2.2791592e-11 * 6.4268857e-24 = 3546288500000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000010100010010110000100110100;
		b = 32'b10011000101000100101100100110010;
		correct = 32'b01101001010110001010000011000000;
		#400 //-68.68985 * -4.1966083e-24 = 1.6367944e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010111011010110110110111000010;
		b = 32'b01000001111000100000010100111000;
		correct = 32'b00010101000001010101010000000001;
		#400 //7.607113e-25 * 28.252548 = 2.6925403e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011011101101110100000111111000;
		b = 32'b11010100000100100111000111000110;
		correct = 32'b11000111001000000010110100111100;
		#400 //1.0316491e+17 * -2515896000000.0 = -41005.234
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011110000101011100110010011001;
		b = 32'b01100010100011111100110111010101;
		correct = 32'b10111011000001010101011000011000;
		#400 //-2.6985427e+18 * 1.3263581e+21 = -0.0020345505
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010010001110001100001111111100;
		b = 32'b10010100011000000010100011110111;
		correct = 32'b11111101010100110000001010001001;
		#400 //198390510000.0 * -1.1317189e-26 = -1.7530017e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110001110101010101100111111100;
		b = 32'b11100100001100000100001100111000;
		correct = 32'b10001101000110101110111011111111;
		#400 //6.209346e-09 * -1.3005882e+22 = -4.7742595e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010000100000110100010000011011;
		b = 32'b00110111110001011100101111011101;
		correct = 32'b01011000001010011110010001111000;
		#400 //17618230000.0 * 2.3579161e-05 = 747194900000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011010101111110111000100000110;
		b = 32'b01010101100110110101000111010111;
		correct = 32'b10000100100111011100010010101011;
		#400 //-7.917835e-23 * 21346975000000.0 = -3.7091134e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011001100000100110111010000101;
		b = 32'b01010110101000010011100110110101;
		correct = 32'b01000010010011110001101011000101;
		#400 //4589158000000000.0 * 88634610000000.0 = 51.776142
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001110110101110010111110000101;
		b = 32'b10111100111001101110111110111010;
		correct = 32'b01010001011011101000101000101101;
		#400 //-1805107800.0 * -0.028190482 = 64032526000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100100010000111111001111110000;
		b = 32'b00101011100111001101101011111111;
		correct = 32'b00111000000111111110011110101101;
		#400 //4.2490508e-17 * 1.114525e-12 = 3.812432e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111101111010000101001101000011;
		b = 32'b11001001101001100010010011100000;
		correct = 32'b01110011101100101111110010101111;
		#400 //-3.8601652e+37 * -1361052.0 = 2.836163e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000011001001000111101000101000;
		b = 32'b11000000001111101011110000010100;
		correct = 32'b00000010010111001100000111111011;
		#400 //-4.8335497e-37 * -2.9802294 = 1.6218717e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101011111100010011010100000111;
		b = 32'b00110011110111000000000101101110;
		correct = 32'b00110111100011000101010111001011;
		#400 //1.7138798e-12 * 1.02448084e-07 = 1.6729251e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001010010000011001001101011110;
		b = 32'b10111111111001000111000011000011;
		correct = 32'b01001001110110001110110111010100;
		#400 //-3171543.5 * -1.7846912 = 1777082.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011110101101001100110010010011;
		b = 32'b01001011111000010011111100110000;
		correct = 32'b00010010010011010111101111011010;
		#400 //1.9142851e-20 * 29523552.0 = 6.4839253e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100101101100100110100001101011;
		b = 32'b10000101011001111000111100010110;
		correct = 32'b11011111110001010011110100100110;
		#400 //3.0948834e-16 * -1.08878485e-35 = -2.8425116e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110011001111010011010101001;
		b = 32'b11100111110000111110101011100110;
		correct = 32'b10010110000101110101100010010000;
		#400 //0.2262217 * -1.8503892e+24 = -1.2225628e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011010011110110001111011111111;
		b = 32'b10101000110101011100110010100100;
		correct = 32'b00110001000101100101100000011110;
		#400 //-5.1930622e-23 * -2.3736499e-14 = 2.1877962e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100001111101100101100110011001;
		b = 32'b00110000001000101001011000110010;
		correct = 32'b11110001010000011111000111001100;
		#400 //-5.680444e+20 * 5.9148697e-10 = -9.6036674e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011111010001000101011010000110;
		b = 32'b10110110000101011111111110110000;
		correct = 32'b01101000101001111000101100001001;
		#400 //-1.4147643e+19 * -2.235156e-06 = 6.3295996e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101100101110101100110110011111;
		b = 32'b00011010111101000111110100011111;
		correct = 32'b11010001010000111001100100110100;
		#400 //-5.3092665e-12 * 1.0111818e-22 = -52505560000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110101010000111000011001001000;
		b = 32'b11010110010111101101110101101000;
		correct = 32'b10011110011000001001100001000010;
		#400 //7.2838566e-07 * -61260630000000.0 = -1.18899474e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010000110111010010101000011011;
		b = 32'b10000101000001001010110000101101;
		correct = 32'b11001011010101010110000000010110;
		#400 //8.7234004e-29 * -6.238234e-36 = -13983766.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011111000111111000100110100111;
		b = 32'b11000001010000100011111111000100;
		correct = 32'b11011101010100100100000100001000;
		#400 //1.1495903e+19 * -12.140568 = -9.4689996e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110001010110100110000000111010;
		b = 32'b00010001111111101010100000100100;
		correct = 32'b11011110110110111000011100011001;
		#400 //-3.1777874e-09 * 4.0177759e-28 = -7.90932e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001000010001111011010000101101;
		b = 32'b00110010110011011100110010001110;
		correct = 32'b01010100111110000110101011111111;
		#400 //204496.7 * 2.3958162e-08 = 8535576000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010100101110100001110111111111;
		b = 32'b11010011000010011000001010011111;
		correct = 32'b10000001001011010011111011001010;
		#400 //1.8793032e-26 * -590602000000.0 = -3.182013e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011100110000111111010001101111;
		b = 32'b11000101100100001101000110100100;
		correct = 32'b10010110101011010011001001110110;
		#400 //1.2967202e-21 * -4634.205 = -2.7981503e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001000111011001001110000010000;
		b = 32'b10110110000101000101011111001010;
		correct = 32'b11010010010011000010100110001100;
		#400 //484576.5 * -2.2104819e-06 = -219217600000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000101010110011101010110101010;
		b = 32'b10111001011011101111010101011000;
		correct = 32'b01001011011010010101111010101010;
		#400 //-3485.354 * -0.00022788846 = 15294122.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001101111110111101110111001110;
		b = 32'b01000010111110110011110100011100;
		correct = 32'b01001010100000000101000111011111;
		#400 //528202180.0 * 125.619354 = 4204783.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100111010011010001001011111010;
		b = 32'b11101010110100001011001011110101;
		correct = 32'b10111011111110111000110110110010;
		#400 //9.684352e+23 * -1.2615084e+26 = -0.0076768035
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001100000000111110101110011011;
		b = 32'b01001010110011010101101011000010;
		correct = 32'b01000000101001000111010010000100;
		#400 //34582124.0 * 6729057.0 = 5.139223
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110101100010011110010010000101;
		b = 32'b11100100010110011010000010100111;
		correct = 32'b01010000101000100011010011000100;
		#400 //-3.495994e+32 * -1.6058079e+22 = 21770936000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000000011100010000111110010111;
		b = 32'b10001100101100110001100111010111;
		correct = 32'b10110011001000011001101011011011;
		#400 //1.0383004e-38 * -2.7594869e-31 = -3.7626574e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011010111110101011000110111101;
		b = 32'b01000101011011001000011111101010;
		correct = 32'b10010101000001111010101000100010;
		#400 //-1.0368473e-22 * 3784.4946 = -2.7397244e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011000100100010011110011101110;
		b = 32'b10100001111001111110011001011011;
		correct = 32'b10110110001000000101010011110101;
		#400 //3.7543145e-24 * -1.5714143e-18 = -2.389131e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011000011000001100111000011010;
		b = 32'b00010111101011011100101010101110;
		correct = 32'b11000000001001011001001001110010;
		#400 //-2.9055376e-24 * 1.1231027e-24 = -2.5870633
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100100000001101111100011110101;
		b = 32'b00101000101110110000100001001111;
		correct = 32'b00111010101110001011111000111100;
		#400 //2.9267493e-17 * 2.0764774e-14 = 0.001409478
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011100001110111101010111110010;
		b = 32'b01111101011100111011111110010111;
		correct = 32'b00011110010001010100011011100111;
		#400 //2.1148422e+17 * 2.0249825e+37 = 1.04437554e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100101000100101110011010001011;
		b = 32'b01001111001101001110101000101110;
		correct = 32'b11010101010011111101111001101101;
		#400 //-4.335739e+22 * 3035246000.0 = -14284639000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111101110001011101000000011010;
		b = 32'b01000111011001110011001111011001;
		correct = 32'b11110101110110110000011101111001;
		#400 //-3.2867305e+37 * 59187.848 = -5.5530497e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010000100100010110110101101011;
		b = 32'b10110101010000010100001110110000;
		correct = 32'b11011010110000001010001001110111;
		#400 //19518937000.0 * -7.19966e-07 = -2.7110914e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011000111100000101101000011011;
		b = 32'b11011100001000000101110100110000;
		correct = 32'b10111100001111111101100001011001;
		#400 //2114158300000000.0 * -1.8055383e+17 = -0.011709296
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111000011110010010001001001001;
		b = 32'b00010101010010100110100100000000;
		correct = 32'b01100010100111011000110000010010;
		#400 //5.9398157e-05 * 4.0876406e-26 = 1.453116e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011100001011100011110010001000;
		b = 32'b00110100001101110110011100101000;
		correct = 32'b10100111011100110011010010000001;
		#400 //-5.7650005e-22 * 1.7080731e-07 = -3.3751487e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010010111000011110011100100100;
		b = 32'b00110111001010101010010010100001;
		correct = 32'b10011011001010010111001101011010;
		#400 //-1.4256477e-27 * 1.017112e-05 = -1.4016624e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111100010111101111000011101100;
		b = 32'b11111000011101110101011010010011;
		correct = 32'b10000011011001101011111110100000;
		#400 //0.013607245 * -2.0066457e+34 = -6.78109e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000001011100101000101101100100;
		b = 32'b11000011001101100001001101101010;
		correct = 32'b00111101101010101000001001111011;
		#400 //-15.159031 * -182.07584 = 0.083256684
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101110110000110101011010001100;
		b = 32'b00111101001111100011010010011000;
		correct = 32'b11110001000000110111010000111100;
		#400 //-3.0227103e+28 * 0.046436876 = -6.509289e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101001101111111000000110101111;
		b = 32'b11100010010000011010100110111000;
		correct = 32'b01000110111111010010011001000110;
		#400 //-2.8939656e+25 * -8.931128e+20 = 32403.137
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111111011100010001111010001;
		b = 32'b10000110010100010000110010010111;
		correct = 32'b01110001000100011100111111101000;
		#400 //-2.838849e-05 * -3.931778e-35 = 7.220267e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011111000100111111111100010110;
		b = 32'b10111100010101000101110100100010;
		correct = 32'b11100010001100100110100000010010;
		#400 //1.0664267e+19 * -0.012961658 = -8.227549e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111000101110101000001011111000;
		b = 32'b11111001001001100101000001110011;
		correct = 32'b10111111000011111000101101100000;
		#400 //3.0263237e+34 * -5.397206e+34 = -0.56072044
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100010111000011010011000100000;
		b = 32'b11010001111100101100111000010110;
		correct = 32'b10010000011011011110100101011101;
		#400 //6.1162264e-18 * -130354954000.0 = -4.6919785e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000101101111110110010011010001;
		b = 32'b11010100001101111010111101111010;
		correct = 32'b00110001000001010101111100011100;
		#400 //-6124.602 * -3155692000000.0 = 1.940811e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111110000101001110100101010100;
		b = 32'b01001111101111110011011001000000;
		correct = 32'b11101101110001110101110111101110;
		#400 //-4.9484313e+37 * 6416007000.0 = -7.712634e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101001101101110011010100100101;
		b = 32'b11011100101100000110011111111011;
		correct = 32'b11001100100001001110111101100011;
		#400 //2.768555e+25 * -3.972314e+17 = -69696280.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011000000011100001100011001101;
		b = 32'b11010101011000001100100001010101;
		correct = 32'b00000010001000011101010011000001;
		#400 //-1.8365591e-24 * -15446939000000.0 = 1.1889469e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111011010001100000001010011001;
		b = 32'b01110110010011100100000111011100;
		correct = 32'b11000100011101011100001110010010;
		#400 //-1.0281275e+36 * 1.0458486e+33 = -983.0558
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110010000110111000110001101100;
		b = 32'b01100110011110111010100100100011;
		correct = 32'b10001011000111100011101100001001;
		#400 //-9.054116e-09 * 2.971085e+23 = -3.0474106e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101100110001110101010001010110;
		b = 32'b01010010011011011010010011001101;
		correct = 32'b00011001110101101011100111100111;
		#400 //5.6652833e-12 * 255168040000.0 = 2.2202167e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101100011110000010011101101111;
		b = 32'b11001010001110110101100011101110;
		correct = 32'b00100001101010011000101101100100;
		#400 //-3.526481e-12 * -3069499.5 = 1.1488782e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101111010001000010000011010011;
		b = 32'b11001000011111010111111100101010;
		correct = 32'b10100110010001100001000010100010;
		#400 //1.7837758e-10 * -259580.66 = -6.871759e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110011110110111110010101001111;
		b = 32'b11111010000010110110101011110001;
		correct = 32'b10111001010010011110001100011110;
		#400 //3.484387e+31 * -1.8097457e+35 = -0.00019253462
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001100010011001111011100110110;
		b = 32'b10110111011100111011000000010010;
		correct = 32'b01010100010101110101001001001100;
		#400 //-53730520.0 * -1.4524923e-05 = 3699194700000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101011011110010000001011001000;
		b = 32'b10110001110101111100001100110010;
		correct = 32'b00111001000100111011100101110101;
		#400 //-8.846643e-13 * -6.2795147e-09 = 0.000140881
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110011000011011100111010000110;
		b = 32'b11010110111101010010000100110000;
		correct = 32'b10011011100101000001100001011111;
		#400 //3.3016953e-08 * -134761440000000.0 = -2.4500296e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101000100011000010111100111101;
		b = 32'b01000100010001100101110011101010;
		correct = 32'b11100011101101001110101011000100;
		#400 //-5.2960216e+24 * 793.4518 = -6.674661e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110111101100011001011010010;
		b = 32'b01001010101001001101000000110011;
		correct = 32'b00110011101111110011010011101101;
		#400 //0.48085648 * 5400601.5 = 8.903758e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011011011011111010100101100101;
		b = 32'b10001011111101001100111100100001;
		correct = 32'b01001110111110101001111000000111;
		#400 //-1.9824351e-22 * -9.4297034e-32 = 2102330200.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100100011111001000000111110;
		b = 32'b00100111101101101011001100000111;
		correct = 32'b01011100010010010010100110010110;
		#400 //1148.5076 * 5.070925e-15 = 2.2648878e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100110010001100100110111101011;
		b = 32'b11001010100101110110111010010111;
		correct = 32'b00011011001001111001111010011001;
		#400 //-6.880065e-16 * -4962123.5 = 1.3865162e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010100000010000101001000010001;
		b = 32'b00010111011111111001101011001010;
		correct = 32'b10111100000010001000100000001011;
		#400 //-6.88243e-27 * 8.2590315e-25 = -0.008333216
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000101010101001011010110011;
		b = 32'b00011011000101101100101010011100;
		correct = 32'b11010101000100001100111000010010;
		#400 //-1.2411959e-09 * 1.2473176e-22 = -9950921000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101000001111011010100100001001;
		b = 32'b00011001000110000010000011001001;
		correct = 32'b01001110100111111001010001011001;
		#400 //1.0528261e-14 * 7.864837e-24 = 1338649700.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010011100100010110100000011110;
		b = 32'b11101100101001100111110011010001;
		correct = 32'b00100110010111111001010111000001;
		#400 //-1249034100000.0 * -1.6101689e+27 = 7.757162e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011011110111101010011010010001;
		b = 32'b10011100101110001001001100011001;
		correct = 32'b11111110100110100110011110111101;
		#400 //1.2534117e+17 * -1.2214122e-21 = -1.0261988e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011100110011111010110010010100;
		b = 32'b00101010100000101001110001010101;
		correct = 32'b11110001110010111000010111101010;
		#400 //-4.6764057e+17 * 2.3201116e-13 = -2.0155952e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101101110001111001110001100000;
		b = 32'b00110001110100010010001111000010;
		correct = 32'b11111011011101000101011000001011;
		#400 //-7.7220703e+27 * 6.0867658e-09 = -1.2686656e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010111111001111010111111100000;
		b = 32'b01101111110011010011111001010000;
		correct = 32'b00100111100100000111110111010110;
		#400 //509485130000000.0 * 1.2703952e+29 = 4.010446e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110100000000011100101101010011;
		b = 32'b01001101110010000001000000110100;
		correct = 32'b11100101101001100001010110000101;
		#400 //-4.1133435e+31 * 419563140.0 = -9.8038725e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100100100101011011111001001101;
		b = 32'b10010110010001001010000000101101;
		correct = 32'b01001101110000101111010111110111;
		#400 //-6.494083e-17 * -1.5883296e-25 = 408862430.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000001010010011000010011111101;
		b = 32'b11101111101010011110110000100011;
		correct = 32'b00010001000101111100110100110110;
		#400 //-12.594968 * -1.0517688e+29 = 1.1975035e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100100101001001101100011111110;
		b = 32'b11100011011101011000000000111011;
		correct = 32'b01000000101010111110010111000011;
		#400 //-2.4327216e+22 * -4.5286923e+21 = 5.371797
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101010110101001000001010010110;
		b = 32'b11110111100101111011010010010011;
		correct = 32'b00110010101100110100110110101110;
		#400 //-1.2845447e+26 * -6.153901e+33 = 2.0873667e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001011101000111110000101011101;
		b = 32'b00001111000011100101010001101101;
		correct = 32'b10111100000100110110000101111110;
		#400 //-6.3124405e-32 * 7.0174e-30 = -0.008995412
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000111111111001001011101011101;
		b = 32'b00010000111000011000010101101001;
		correct = 32'b00110110100011110101110101000011;
		#400 //3.800571e-34 * 8.89524e-29 = 4.272589e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110011100101101010100100000010;
		b = 32'b10110100011011110110111101101101;
		correct = 32'b00111110101000010001010101001111;
		#400 //-7.015662e-08 * -2.2299146e-07 = 0.3146157
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011010010000100111101000101;
		b = 32'b11100000000101101110011111000001;
		correct = 32'b00101010101010011110011111001101;
		#400 //-13127493.0 * -4.349549e+19 = 3.0181275e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100010100010101110011101000001;
		b = 32'b10101010011001111111010100100100;
		correct = 32'b11110111100110010100110011111001;
		#400 //1.2811571e+21 * -2.0601972e-13 = -6.218614e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011000100000001010100001010;
		b = 32'b11010100110010110110011111000001;
		correct = 32'b00110101101101010101011001110001;
		#400 //-9442570.0 * -6988952500000.0 = 1.3510709e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000110010101101100100110111011;
		b = 32'b10110010110000111100101101111101;
		correct = 32'b00010011000011000110101010101011;
		#400 //-4.0397135e-35 * -2.2793524e-08 = 1.7723076e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101001000011000100011101111010;
		b = 32'b00111010011101001100010000101011;
		correct = 32'b00101110000100101011011110101001;
		#400 //3.114824e-14 * 0.00093370926 = 3.335968e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111101011110110000010100001100;
		b = 32'b11110110101101111110011001000110;
		correct = 32'b00000110001011101011011111000100;
		#400 //-0.06128411 * -1.8649625e+33 = 3.2860772e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110000110011110011000101111000;
		b = 32'b11011110111000010111000000011011;
		correct = 32'b11010001011010110100100000101101;
		#400 //5.129856e+29 * -8.122257e+18 = -63158014000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001101111011111111100110110001;
		b = 32'b01011010101001011001111010110111;
		correct = 32'b10110010101110010111011101000000;
		#400 //-503264800.0 * 2.330894e+16 = -2.1591063e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001101000101000000011100000101;
		b = 32'b10110000000011111101100001001010;
		correct = 32'b01011100100000111011100011001001;
		#400 //-155218000.0 * -5.233046e-10 = 2.9661116e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100001001011010001110100000001;
		b = 32'b00110011111111011010000100000101;
		correct = 32'b10101100101011101011101101001100;
		#400 //-5.8653066e-19 * 1.181052e-07 = -4.9661716e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101000101100010110110111110001;
		b = 32'b01010101000001100010011100011011;
		correct = 32'b00010011001010010100101010111000;
		#400 //1.9698627e-14 * 9218907000000.0 = 2.1367638e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000011101010111111110010100001;
		b = 32'b00101110011101111111100011010101;
		correct = 32'b11010100101100011000111000001010;
		#400 //-343.97366 * 5.6382305e-11 = -6100738000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011111000011001000111111100100;
		b = 32'b00001100001111100110010110100111;
		correct = 32'b11010010001111001111111001110010;
		#400 //-2.9765177e-20 * 1.4667657e-31 = -202930680000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111000101110100100111001000101;
		b = 32'b11011011101110101000101011111000;
		correct = 32'b11011100011111111010110010110011;
		#400 //3.0229835e+34 * -1.0501429e+17 = -2.8786402e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111011111011111101011110110000;
		b = 32'b11101110011011001001111100000110;
		correct = 32'b00001101000000011011111000011010;
		#400 //-0.007319413 * -1.8307677e+28 = 3.998002e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010001101101010010010100101001;
		b = 32'b01010101010101111101011011001001;
		correct = 32'b00111011110101101101100111000111;
		#400 //97251566000.0 * 14832343000000.0 = 0.006556723
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011101011001101111101100100101;
		b = 32'b11000011011111101001101000001100;
		correct = 32'b10011001011010000011111111100011;
		#400 //3.0570085e-21 * -254.60175 = -1.2007021e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101110001100101100010100101000;
		b = 32'b10011010110000111100000010111111;
		correct = 32'b11010010111010011100101001011001;
		#400 //4.0647624e-11 * -8.096151e-23 = -502061100000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000011101010100111110111001000;
		b = 32'b10111001010000110100000010111000;
		correct = 32'b11001001110111111000100011100011;
		#400 //340.98267 * -0.00018620759 = -1831196.4
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001011011111010101111001000110;
		b = 32'b10101000110111010010010110011100;
		correct = 32'b11100010000100101010011001010101;
		#400 //16604742.0 * -2.455224e-14 = -6.763025e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111000010111011111000001000100;
		b = 32'b11110111001101101101110100110010;
		correct = 32'b11000000100110110101100111100011;
		#400 //1.8005793e+34 * -3.7089234e+33 = -4.8547225
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011100000101110001000100000011;
		b = 32'b01011100110011001100010100101111;
		correct = 32'b10111110101111001101110001001010;
		#400 //-1.700857e+17 * 4.611016e+17 = -0.36886817
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010111010110000101110100110110;
		b = 32'b11111111111100001010110110101001;
		correct = 32'b11111111111100001010110110101001;
		#400 //-6.9911013e-25 * nan = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011111000111011100000000011111;
		b = 32'b11010100010100111111001110101001;
		correct = 32'b00001010001111101000100011010010;
		#400 //-3.3404962e-20 * -3641304200000.0 = 9.1739e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111001000011010011101111001000;
		b = 32'b10010100010010000111100110001010;
		correct = 32'b11100100001101000101100111001101;
		#400 //0.00013469078 * -1.0121389e-26 = -1.3307539e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001001100101010101010111011000;
		b = 32'b10101011010000101101110100101101;
		correct = 32'b11011101110001000010111111110110;
		#400 //1223355.0 * -6.922959e-13 = -1.7670985e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001100010011001111111111010100;
		b = 32'b00011001000110101111011101000110;
		correct = 32'b11110010101010010101001110110111;
		#400 //-53739344.0 * 8.01155e-24 = -6.707734e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101011100001100110100010000000;
		b = 32'b01011010001100101011111011000010;
		correct = 32'b11010000110000001000000000010110;
		#400 //-3.249791e+26 * 1.2578072e+16 = -25836958000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010000110001010100011110110010;
		b = 32'b10101010101000010000101110001100;
		correct = 32'b11100101100111001100110011000011;
		#400 //26478481000.0 * -2.8607357e-13 = -9.2558295e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110010000111110010101001110010;
		b = 32'b01010010001000111011001001011000;
		correct = 32'b00011111011110001110101000010010;
		#400 //9.264669e-09 * 175767950000.0 = 5.270966e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001110101111110000110000100101;
		b = 32'b10111011011011101101001100011001;
		correct = 32'b01010010110011001100100101110001;
		#400 //-1602622100.0 * -0.0036441742 = 439776480000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010010111010111001101010001000;
		b = 32'b10100110100000101111000011101100;
		correct = 32'b01101011111001100100111111001011;
		#400 //-505954960000.0 * -9.085864e-16 = 5.568595e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111000100101100100111100001101;
		b = 32'b10000000111010100001110101110100;
		correct = 32'b01110111001001000101110000001101;
		#400 //-7.167282e-05 * -2.1500072e-38 = 3.3336082e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010001100101111011100011100111;
		b = 32'b10010100110010010010101011111011;
		correct = 32'b10111100010000010001001110111001;
		#400 //2.3937554e-28 * -2.0312766e-26 = -0.011784487
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100101100111110111111001100111;
		b = 32'b01100001011010010100011010100100;
		correct = 32'b00000011101011110000011111001110;
		#400 //2.7667757e-16 * 2.6894885e+20 = 1.0287367e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110011011010000000101000001001;
		b = 32'b00001001001101011110110011000100;
		correct = 32'b01101001101000110100001010000010;
		#400 //5.4025836e-08 * 2.189841e-33 = 2.4671123e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111011110000011000111010100111;
		b = 32'b10101011111010100101110011100011;
		correct = 32'b11001111010100110110110101010110;
		#400 //0.005906898 * -1.6652481e-12 = -3547158000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000100000101101100001110110110;
		b = 32'b11000000101111000111110000000100;
		correct = 32'b01000010110011001100010011001001;
		#400 //-603.058 * -5.8901386 = 102.384346
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100010101011111010000010011010;
		b = 32'b00010010001001101001101010110110;
		correct = 32'b11010000000001101110111010101001;
		#400 //-4.760389e-18 * 5.257106e-28 = -9055151000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010001011010100101000101111100;
		b = 32'b00010110000001001100110010011010;
		correct = 32'b00111010111000011101100110101100;
		#400 //1.8484454e-28 * 1.0727436e-25 = 0.0017231009
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010000100011001010011101101111;
		b = 32'b10110010101011100001001100110010;
		correct = 32'b10011101010011101101100110100010;
		#400 //5.5478236e-29 * -2.0264995e-08 = -2.7376387e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010001110010111001110011000000;
		b = 32'b01001001110001111100111100110011;
		correct = 32'b01000111100000100110111110101011;
		#400 //109313520000.0 * 1636838.4 = 66783.336
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001101100001111110011000010010;
		b = 32'b11011011010111011110010000111001;
		correct = 32'b10110001100111001100100111100110;
		#400 //285000260.0 * -6.2456903e+16 = -4.5631507e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000100011100100100100101010;
		b = 32'b11001001010000101010100110111001;
		correct = 32'b00100110101110110001111001111110;
		#400 //-1.0352654e-09 * -797339.56 = 1.2983997e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001010111011101110111010101100;
		b = 32'b00001000011110000110011110011011;
		correct = 32'b11000001111101100011110011101100;
		#400 //-2.3008345e-32 * 7.4751573e-34 = -30.779747
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011101111001010100011011111011;
		b = 32'b11010101100011100001011110010010;
		correct = 32'b01000111110011101000100111011110;
		#400 //-2.065146e+18 * -19528986000000.0 = 105747.734
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111011110011000010100011000100;
		b = 32'b10010100001000000110001000100101;
		correct = 32'b01100111001000101110111111011110;
		#400 //-0.0062304456 * -8.097291e-27 = 7.6944814e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101100111000110111101111010100;
		b = 32'b11001110101111011001100110110000;
		correct = 32'b01011101100110011001001101000010;
		#400 //-2.2000874e+27 * -1590483000.0 = 1.3832827e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110010000100010100100100010110;
		b = 32'b00100001101111111110100010111010;
		correct = 32'b01001111110000011100111001000110;
		#400 //8.456729e-09 * 1.3004266e-18 = 6503042000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100110011001111101011111001110;
		b = 32'b01000111100000011100010101001011;
		correct = 32'b01011110011001001010110111111000;
		#400 //2.7371189e+23 * 66442.586 = 4.1195248e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110111100011011101011010101101;
		b = 32'b00011101110100101111010011110111;
		correct = 32'b01011001001011000001111110101001;
		#400 //1.6908476e-05 * 5.5839825e-21 = 3028031700000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010111110011000100011110011000;
		b = 32'b01111111001010010010111100100110;
		correct = 32'b10011000000110101000110101100001;
		#400 //-449215730000000.0 * 2.2488434e+38 = -1.9975412e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000101110100010011011010110001;
		b = 32'b00001000101011011000110100101101;
		correct = 32'b01111100100110100100110101010011;
		#400 //6694.8364 * 1.0445249e-33 = 6.409456e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111100010001111100000000111110;
		b = 32'b01110001001110101110101001011101;
		correct = 32'b10001010100010001100101000101101;
		#400 //-0.01219183 * 9.255606e+29 = -1.3172374e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100100100010000101111001010001;
		b = 32'b01010001011001010100111010010011;
		correct = 32'b00010010100110000011111000100100;
		#400 //5.9140376e-17 * 61554110000.0 = 9.607867e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001110010101000010100101111111;
		b = 32'b10111011111011001110110010010101;
		correct = 32'b00010001111001010011111010000110;
		#400 //-2.6150997e-30 * -0.007230351 = 3.6168363e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011011000010010101000001000001;
		b = 32'b10101101000011101011011000111101;
		correct = 32'b01101101011101100101000011110111;
		#400 //-3.865031e+16 * -8.1122305e-12 = 4.7644496e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010101110100010010000010100001;
		b = 32'b01011111100110011010010101111001;
		correct = 32'b00110101101011100011100001100100;
		#400 //28742259000000.0 * 2.2142777e+19 = 1.2980422e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100101101110100111000101010111;
		b = 32'b01000110010011110011110100010100;
		correct = 32'b11011110111001100100111110100010;
		#400 //-1.10056365e+23 * 13263.27 = -8.2978306e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001010111001111111000111110001;
		b = 32'b10111000011101101000111011111001;
		correct = 32'b00010001111100001101001110110110;
		#400 //-2.2335499e-32 * -5.8784124e-05 = 3.79958e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011100110101001110001000010000;
		b = 32'b01001111011111100111100011001111;
		correct = 32'b01001100110101100010100101010010;
		#400 //4.7937003e+17 * 4269330200.0 = 112282260.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100100101011110110110010000010;
		b = 32'b11000110000101100101011111101101;
		correct = 32'b11011110000101010101101001100001;
		#400 //2.5887992e+22 * -9621.981 = -2.6905052e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110000010110001000011110100;
		b = 32'b10001000101000111101111010001001;
		correct = 32'b01101100110110010100000010001101;
		#400 //-2.0722482e-06 * -9.862523e-34 = 2.1011339e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111000110111101010000001101001;
		b = 32'b01010111011000010001000110011101;
		correct = 32'b11100000111111010011100011100000;
		#400 //-3.6123231e+34 * 247465760000000.0 = -1.4597264e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010111111001100000110001101001;
		b = 32'b00011110000111011000110100001011;
		correct = 32'b01111001001110101110011001001010;
		#400 //505881950000000.0 * 8.340678e-21 = 6.0652377e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100110001101010101100010000101;
		b = 32'b10111001011011011110001101101010;
		correct = 32'b00101100010000110010011100001111;
		#400 //-6.2916956e-16 * -0.000226868 = 2.7732849e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100010111111000011101000001101;
		b = 32'b00101110111001000111001101110011;
		correct = 32'b01110011100011010101001001001011;
		#400 //2.3263813e+21 * 1.03887475e-10 = 2.2393279e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011101101100011110111011110111;
		b = 32'b11010011001011101101010010000010;
		correct = 32'b10001010000000100100010110100111;
		#400 //4.7098594e-21 * -750889600000.0 = -6.2723725e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101110001101001111011111010011;
		b = 32'b11100010001001001110111001000110;
		correct = 32'b01001011100011000111001001000000;
		#400 //-1.4001726e+28 * -7.6060886e+20 = 18408576.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000000000100101011101111100011;
		b = 32'b00111100010101000111110111000011;
		correct = 32'b11000011001100001100011101001100;
		#400 //-2.2927177 * 0.012969437 = -176.7785
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001101001011110110100111111110;
		b = 32'b11001010101010010100111011100010;
		correct = 32'b10000010000001001001110110111101;
		#400 //5.405362e-31 * -5547889.0 = -9.743097e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101101011110100001010011110000;
		b = 32'b11011011000000101011110111010011;
		correct = 32'b01010001111101001101011001111110;
		#400 //-4.8372853e+27 * -3.680046e+16 = 131446325000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001011100100110010100001011111;
		b = 32'b00001110000010100001011111000000;
		correct = 32'b00111101000010000110011100000100;
		#400 //5.6683084e-32 * 1.7021248e-30 = 0.03330137
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011111011011101111011011100111;
		b = 32'b11000000011110001110000101001101;
		correct = 32'b01011110011101011100110011111100;
		#400 //-1.7219204e+19 * -3.8887513 = 4.427952e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110000010101101100000010111011;
		b = 32'b01111101111111101110111010010000;
		correct = 32'b00110001110101111010011100010011;
		#400 //2.6585116e+29 * 4.2357825e+37 = 6.2763177e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110000010000011100100101011111;
		b = 32'b01000100001100110000010100001111;
		correct = 32'b11101011100010101000111011110001;
		#400 //-2.398962e+29 * 716.07904 = -3.3501357e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101011111110001010001010010110;
		b = 32'b10100010000100110101010000111100;
		correct = 32'b01001001010110000000001111011100;
		#400 //-1.7666587e-12 * -1.9966808e-18 = 884797.75
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001111011011001011100010011100;
		b = 32'b10011010100100010011100000110010;
		correct = 32'b00110100010100001010011011011001;
		#400 //-1.1671253e-29 * -6.006138e-23 = 1.9432208e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110000101110001100001011011000;
		b = 32'b11000011000100100100001110100100;
		correct = 32'b10101101001000011011000010010010;
		#400 //1.344314e-09 * -146.26422 = -9.190997e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100010110110100110111001001000;
		b = 32'b10010011111101000000111010011100;
		correct = 32'b11001110011001010001111010100100;
		#400 //5.9205783e-18 * -6.1608665e-27 = -960997600.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000100101011110010101000101001;
		b = 32'b00010010111111110100110110010110;
		correct = 32'b10110001001011111010010010010010;
		#400 //-4.118102e-36 * 1.6111889e-27 = -2.55594e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101010100101000010111000011011;
		b = 32'b00000100101100001011010110011101;
		correct = 32'b11100101010101101010101101011101;
		#400 //-2.6322073e-13 * 4.1544187e-36 = -6.335922e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000111001110100010010101110010;
		b = 32'b01111111110100111000110101100001;
		correct = 32'b01111111110100111000110101100001;
		#400 //-47653.445 * nan = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010100110110011101111000111011;
		b = 32'b11000101000100010110101010110111;
		correct = 32'b01001111001111111100011000001011;
		#400 //-7485890500000.0 * -2326.6697 = 3217427200.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011111101001100001010110111001;
		b = 32'b00011000010000000011101110111010;
		correct = 32'b01000110110111010010110101111110;
		#400 //7.033967e-20 * 2.4845573e-24 = 28310.746
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011000111000011011000000101001;
		b = 32'b00100000111100010100000010001101;
		correct = 32'b01110111011011110111110000001011;
		#400 //1985173700000000.0 * 4.0869704e-19 = 4.8573236e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111110000110010110010010101111;
		b = 32'b00110001011001110010001110100001;
		correct = 32'b11001100001010011110010001010110;
		#400 //-0.14979814 * 3.3635177e-09 = -44536150.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010111110110010111010001110100;
		b = 32'b10100110100000110000000111001001;
		correct = 32'b11110000110101000111011010110101;
		#400 //478188370000000.0 * -9.090435e-16 = -5.2603464e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111011000101001111101001110000;
		b = 32'b00100000001000110110110111101111;
		correct = 32'b01011010011010010101110100000100;
		#400 //0.002273228 * 1.3843011e-19 = 1.6421485e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010010001010111001111101000101;
		b = 32'b00101101100101111101111001000101;
		correct = 32'b00100100000100001010011000111001;
		#400 //5.41544e-28 * 1.726542e-11 = 3.136582e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010110100101010000110000111001;
		b = 32'b11000000101001111101111011110000;
		correct = 32'b10010101011000110100101110001100;
		#400 //2.4079962e-25 * -5.245964 = -4.590188e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001111010000000100001010100100;
		b = 32'b10101000100100110010001111101110;
		correct = 32'b10100110001001110100000000101011;
		#400 //9.4791654e-30 * -1.633586e-14 = -5.802673e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111100010100111011010011100101;
		b = 32'b10110110010001101110111010110000;
		correct = 32'b11000101100010000011100000101010;
		#400 //0.012921547 * -2.9643234e-06 = -4359.0205
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000011101001011000011101001001;
		b = 32'b01110100100101001101111001001010;
		correct = 32'b10001110100011100101001100100001;
		#400 //-331.05692 * 9.435651e+31 = -3.5085753e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011111011111010110100101010001;
		b = 32'b00010001001101100101011110111101;
		correct = 32'b11001101101100011110001101101111;
		#400 //-5.366195e-20 * 1.4384305e-28 = -373059040.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110011010111000001100111011111;
		b = 32'b11100110111011111110110100010100;
		correct = 32'b01001011111010101101100011000111;
		#400 //-1.7438202e+31 * -5.6650945e+23 = 30781838.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110110001010010111110101000;
		b = 32'b11100110011001100001010010111100;
		correct = 32'b00001111110110110110011001000110;
		#400 //-5.8766054e-06 * -2.716317e+23 = 2.1634462e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101111111010011101011001011000;
		b = 32'b01011110111100101001101111100011;
		correct = 32'b00010000011101101011111010000011;
		#400 //4.2534753e-10 * 8.740908e+18 = 4.866171e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101111110001110000101100100110;
		b = 32'b11010011000001010011011111111001;
		correct = 32'b00011100001111110011111100001110;
		#400 //-3.620581e-10 * -572169700000.0 = 6.3278095e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111101111101111110100101110000;
		b = 32'b10001000001111111000001000111101;
		correct = 32'b01110101001001011011001011010011;
		#400 //-0.121050715 * -5.7630066e-34 = 2.1004784e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001100001111011011101101100100;
		b = 32'b10111000100000011110011110000101;
		correct = 32'b10010011001110101111001101011000;
		#400 //1.4616421e-31 * -6.194323e-05 = -2.3596478e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010001010010111011000011101110;
		b = 32'b10111001100000110100010101001001;
		correct = 32'b00010111010001101001110110111001;
		#400 //-1.6068397e-28 * -0.0002503789 = 6.4176324e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010101010010111101101011111011;
		b = 32'b01001000111011000110110110111001;
		correct = 32'b10001011110111001011101011111100;
		#400 //-4.116827e-26 * 484205.78 = -8.502226e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001010111110001111100101111000;
		b = 32'b10110010001001001100001101000101;
		correct = 32'b01011000010000010110110000000100;
		#400 //-8158396.0 * -9.5904555e-09 = 850678700000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101101000111011000001101010000;
		b = 32'b01010110011010001100000101101110;
		correct = 32'b10010110001011010011111001000000;
		#400 //-8.953574e-12 * 63979370000000.0 = -1.3994471e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110001011101101011000000111001;
		b = 32'b11101110000101011100000000010100;
		correct = 32'b01000010110100101101101111000001;
		#400 //-1.22154164e+30 * -1.1586369e+28 = 105.42921
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101011001110111100110100111000;
		b = 32'b01110100100110011101010111010001;
		correct = 32'b10110110000111000100001100010111;
		#400 //-2.2703825e+26 * 9.750465e+31 = -2.3284863e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010000110111001110111001111001;
		b = 32'b00101101110100001111000010110101;
		correct = 32'b01100010100001110101100010010110;
		#400 //29652929000.0 * 2.3753758e-11 = 1.2483469e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111100001110010111010010000000;
		b = 32'b01101111101101001100010100101001;
		correct = 32'b01001100000000110101000100111011;
		#400 //3.8517513e+36 * 1.1189131e+29 = 34424044.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111110101110101011010000110110;
		b = 32'b11000110110010011010110011100010;
		correct = 32'b01110111011011001111111011101111;
		#400 //-1.2408606e+38 * -25814.441 = 4.8068466e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011100110011101011010010000001;
		b = 32'b01000110000001000101111110010111;
		correct = 32'b11010110010001111110000000111011;
		#400 //-4.654585e+17 * 8471.897 = -54941470000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100001101100110001100100110;
		b = 32'b00101011000010010001011010011000;
		correct = 32'b01011000101010100100101111000011;
		#400 //729.5492 * 4.870353e-13 = 1497939000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101111000111100000000111001000;
		b = 32'b01100101111101100110101100011011;
		correct = 32'b10001000101001000010011010011101;
		#400 //-1.4370649e-10 * 1.4545974e+23 = -9.879469e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000000101011001111110000001011;
		b = 32'b10000000000001110111010010110100;
		correct = 32'b11000001101110011001101111100011;
		#400 //1.5886121e-38 * -6.84714e-40 = -23.201117
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111100010001000001110111110111;
		b = 32'b01010111010110000110001100000001;
		correct = 32'b01100100011010000000010100000101;
		#400 //4.0731918e+36 * 237919730000000.0 = 1.7120025e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010010100111111100101011100101;
		b = 32'b10111110010111100101011011011110;
		correct = 32'b01010011101101111111101111101100;
		#400 //-343151900000.0 * -0.21712825 = 1580411100000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110110111100100001111100000100;
		b = 32'b10110100001011000001101101010100;
		correct = 32'b11000010001101000001001001001001;
		#400 //7.2157727e-06 * -1.602869e-07 = -45.017857
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010010110110011011011001011010;
		b = 32'b01001010010010110110110101010010;
		correct = 32'b00001000000010001111110100010010;
		#400 //1.3739578e-27 * 3332948.5 = 4.1223494e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011000111010010100010111101000;
		b = 32'b11001011001111000100110010000111;
		correct = 32'b11001101000111101001001001110100;
		#400 //2051891600000000.0 * -12340359.0 = -166274880.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111011100101010010001100010111;
		b = 32'b00110000011110001011000111110110;
		correct = 32'b01001010100110011000010010000011;
		#400 //0.004551302 * 9.047477e-10 = 5030465.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001001001101000011101010110100;
		b = 32'b10010100000110000001110001011000;
		correct = 32'b00110100100101111010100101011101;
		#400 //-2.1694314e-33 * -7.679629e-27 = 2.824917e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000001111100000101101111101100;
		b = 32'b00000000000001010011011001110010;
		correct = 32'b01000011001110000111000100100011;
		#400 //8.829398e-38 * 4.78709e-40 = 184.44194
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011001100010000010101111110011;
		b = 32'b00111010010110011011110000010011;
		correct = 32'b11011110101000000001101001010111;
		#400 //-4791115000000000.0 * 0.00083059183 = -5.7683145e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111000001001110100000010011111;
		b = 32'b01101000000000100110100010001010;
		correct = 32'b00001111101001000010100111100100;
		#400 //3.9876086e-05 * 2.4633442e+24 = 1.6187784e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100010001111010000101101001110;
		b = 32'b10100110101000100000101001000111;
		correct = 32'b00111011000101010101010011001011;
		#400 //-2.562026e-18 * -1.1243794e-15 = 0.0022786136
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100000110101010000010100100010;
		b = 32'b11100000001010101001011010000000;
		correct = 32'b11000000000111111101011010111101;
		#400 //1.227977e+20 * -4.916861e+19 = -2.4974816
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110101100000010100011101100101;
		b = 32'b00011101001001000011001000100001;
		correct = 32'b01010111110010011000111101111110;
		#400 //9.632028e-07 * 2.1731135e-21 = 443236260000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110111100110000001111010000100;
		b = 32'b10011001110000101100111101000111;
		correct = 32'b11011101010001111110011001111011;
		#400 //1.8134022e-05 * -2.0142849e-23 = -9.00271e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100001011011011101111010001011;
		b = 32'b11011001000100001100110110100100;
		correct = 32'b01000111110100100100010000110110;
		#400 //-2.7424464e+20 * -2547406300000000.0 = 107656.42
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011101010100010000101001000000;
		b = 32'b01100000001101100001011010010110;
		correct = 32'b00111100100100101111001000101001;
		#400 //9.4143264e+17 * 5.248336e+19 = 0.017937737
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101100110110000101000000000001;
		b = 32'b01010001100111100001001001101100;
		correct = 32'b11011010101011110010100100100110;
		#400 //-2.0920463e+27 * 84864240000.0 = -2.4651682e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110101011101010110110001001011;
		b = 32'b11100011000100110111101000111011;
		correct = 32'b00010001110101010000001010000011;
		#400 //-9.14272e-07 * -2.720479e+21 = 3.3607023e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111111010011101110010101101101;
		b = 32'b01110110001000010100101111011100;
		correct = 32'b00001000101001000010111111001100;
		#400 //0.80818826 * 8.178695e+32 = 9.881628e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000011100110111001110010100001;
		b = 32'b00111100100011110010010111100111;
		correct = 32'b00000110100010110010010100010101;
		#400 //9.1460415e-37 * 0.017474128 = 5.2340476e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101001100100011001100111101101;
		b = 32'b01101110110001000110100101000100;
		correct = 32'b10111010001111011100011001100100;
		#400 //-2.2002642e+25 * 3.039316e+28 = -0.00072393403
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000111101110001100110010101111;
		b = 32'b00011010001001110101011100101011;
		correct = 32'b11101101000011010101101011000100;
		#400 //-94617.37 * 3.4605204e-23 = -2.7341947e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100111100010101011100011011111;
		b = 32'b10111001001101101010001001000011;
		correct = 32'b10101101110000100111001011001111;
		#400 //3.850313e-15 * -0.0001741732 = -2.2106232e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000110101001110100101010001011;
		b = 32'b01000011001101101001110111011100;
		correct = 32'b10000010111010101000010000100000;
		#400 //-6.292795e-35 * 182.61664 = -3.4459046e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001001000000100110001100101011;
		b = 32'b00100011100000001001000001110011;
		correct = 32'b11100101000000011101000010101100;
		#400 //-534066.7 * 1.3938964e-17 = -3.831466e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001111100101011000110100110011;
		b = 32'b00111110100000001001001111001111;
		correct = 32'b01010000100101001110000101001000;
		#400 //5018117600.0 * 0.2511277 = 19982336000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101000100101100100111111101000;
		b = 32'b00111011111110000010101100101110;
		correct = 32'b10101100000110110000111000110010;
		#400 //-1.6688e-14 * 0.007573507 = -2.2034705e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010001100100101001000001111110;
		b = 32'b01001011100001011111101010100110;
		correct = 32'b01000101100011000000011000010000;
		#400 //78686175000.0 * 17560908.0 = 4480.758
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010001110110110100111000110100;
		b = 32'b00101110000011011110111100111010;
		correct = 32'b10100011010001011100011001101011;
		#400 //-3.4600304e-28 * 3.2272164e-11 = -1.0721408e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111000010101001111000101001101;
		b = 32'b00100101000110000111000111101101;
		correct = 32'b11010010101100101100101111101101;
		#400 //-5.0769468e-05 * 1.3222498e-16 = -383962740000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111000110100111111100101110011;
		b = 32'b11101111001111101110100000110110;
		correct = 32'b01001001000011100010000000010011;
		#400 //-3.4394815e+34 * -5.908288e+28 = 582145.2
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001111100000100001010010011101;
		b = 32'b00110100011010010010100100111010;
		correct = 32'b11011010100011101101001010000111;
		#400 //-4364778000.0 * 2.1714814e-07 = -2.0100462e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111100010111100001100011100101;
		b = 32'b01000001100001000111011011010100;
		correct = 32'b00111010010101101001110011000011;
		#400 //0.01355574 * 16.558022 = 0.00081868115
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000101011001101111010000001101;
		b = 32'b01100111100001001101110001000100;
		correct = 32'b10011101010111101000000100100000;
		#400 //-3695.2532 * 1.2548311e+24 = -2.9448211e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011111110110111011010010001000;
		b = 32'b00000010100011100010111000001010;
		correct = 32'b01011100110001011100101100101011;
		#400 //9.304877e-20 * 2.089145e-37 = 4.4539165e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111110010001101100101000101010;
		b = 32'b01001111110101101011011010100000;
		correct = 32'b01101101111011010000001110110000;
		#400 //6.605921e+37 * 7204585500.0 = 9.1690507e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100111110010100010001001001100;
		b = 32'b00010010011110100000111011000111;
		correct = 32'b11010100110011101110111111111010;
		#400 //-5.6103447e-15 * 7.8904305e-28 = -7110315000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101100011101010110011011011101;
		b = 32'b01011000101010111010111000100101;
		correct = 32'b10010011001101101111011011111001;
		#400 //-3.4873695e-12 * 1510115500000000.0 = -2.3093396e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011001000100111110011111011100;
		b = 32'b11001101001000010110000011010011;
		correct = 32'b00001011011010101010000011001001;
		#400 //-7.6465455e-24 * -169217330.0 = 4.5187722e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100111100110010001110111011010;
		b = 32'b11111000110010101101011010011111;
		correct = 32'b00101110010000010011111100101010;
		#400 //-1.4461455e+24 * -3.2912406e+34 = 4.393922e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001001111100000100101000110010;
		b = 32'b11010101000010110011101101101011;
		correct = 32'b00110100010111001110011110111100;
		#400 //-1968454.2 * -9567957000000.0 = 2.0573401e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110110000010111110011111010101;
		b = 32'b01101001100101111101010101110000;
		correct = 32'b11001011111010111110001101110100;
		#400 //-7.0940564e+32 * 2.2944466e+25 = -30918376.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101110101001000000011101001001;
		b = 32'b01010001110101010011100100001001;
		correct = 32'b01011100010001001110111110101010;
		#400 //2.5382174e+28 * 114473116000.0 = 2.2173044e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010110111001111101011001101100;
		b = 32'b00110101101011111110001001000111;
		correct = 32'b11100000101010001011100001110000;
		#400 //-127454060000000.0 * 1.3104371e-06 = -9.726072e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111010100001001001101001110101;
		b = 32'b10011100010101100001010111110011;
		correct = 32'b11011101100111101001000010010101;
		#400 //0.0010116833 * -7.083503e-22 = -1.4282245e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010010100000010000111111011011;
		b = 32'b00001111110111100110010111100110;
		correct = 32'b01000010000101001000111111010011;
		#400 //8.144953e-28 * 2.193014e-29 = 37.140453
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100001110011000010010101001000;
		b = 32'b11100000001101110111001011110001;
		correct = 32'b10000001000011100111000011011111;
		#400 //1.3833446e-18 * -5.287557e+19 = -2.6162262e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101010110001010110101001111111;
		b = 32'b01000001010001111110111000110111;
		correct = 32'b10101000111111001100011111000001;
		#400 //-3.5068126e-13 * 12.495658 = -2.806425e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111110011101110111110010111110;
		b = 32'b00100100100101110111001100011110;
		correct = 32'b11011001010100010010101011101010;
		#400 //-0.24168679 * 6.568083e-17 = -3679716000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100011000111100111001110101111;
		b = 32'b11101001110011100111011100111111;
		correct = 32'b10111000110001000111011110000011;
		#400 //2.9229214e+21 * -3.120023e+25 = -9.368269e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100100110100000011100101010001;
		b = 32'b11110000010101110101011100100100;
		correct = 32'b10110011111101111000101000110000;
		#400 //3.0728423e+22 * -2.665785e+29 = -1.152697e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001110010011111110111100001111;
		b = 32'b10011000001101101000100001101011;
		correct = 32'b11110101100100011100111111101111;
		#400 //872137660.0 * -2.3591822e-24 = -3.6967795e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110011101000010100011000001000;
		b = 32'b11010101011100111011101010000001;
		correct = 32'b10011101101010010110010010111101;
		#400 //7.509885e-08 * -16748897000000.0 = -4.483809e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001010111101111110011100000100;
		b = 32'b01111101100011000100100000101100;
		correct = 32'b10001100111000100011001010111000;
		#400 //-8123266.0 * 2.3308332e+37 = -3.4851339e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011100101100001100010011011000;
		b = 32'b11100110110110000000110110000111;
		correct = 32'b00110101010100010111001111100010;
		#400 //-3.9804822e+17 * -5.1014035e+23 = 7.80272e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110111000001010000001011000;
		b = 32'b10100111100110010010111111110100;
		correct = 32'b11010110101110111011000101100010;
		#400 //0.43872333 * -4.251802e-15 = -103185260000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010100100010001011101010100110;
		b = 32'b11100001111100010111000110001101;
		correct = 32'b00110010000100001111100011101110;
		#400 //-4697976000000.0 * -5.5673094e+20 = 8.438503e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101010100000100010100000100011;
		b = 32'b00101110011100010110000100111111;
		correct = 32'b11111011100010100000101001001110;
		#400 //-7.867495e+25 * 5.4883428e-11 = -1.433492e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110011000101011000001111011101;
		b = 32'b00101001000011000100001011101101;
		correct = 32'b11001001100010000111000111011001;
		#400 //-3.4811695e-08 * 3.1144294e-14 = -1117755.1
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000110000111001101000100101110;
		b = 32'b01001101001001110001100010101100;
		correct = 32'b10111000011100000100000001101100;
		#400 //-10036.295 * 175213250.0 = -5.7280457e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111001001011100111011100010001;
		b = 32'b11011111011101100100100110011111;
		correct = 32'b00011001001101010101100001011110;
		#400 //-0.00016638289 * -1.7746891e+19 = 9.375326e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001111000001011010110110101111;
		b = 32'b00111010010010101011111000110100;
		correct = 32'b01010100001010001100101100011110;
		#400 //2242752300.0 * 0.0007734031 = 2899849000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100000101110101111000001100110;
		b = 32'b10110100111110011110111111011111;
		correct = 32'b10101011001111110111100101001110;
		#400 //3.1668708e-19 * -4.6554393e-07 = -6.8025175e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001101011000011111010110000001;
		b = 32'b10111000110001111011000110100101;
		correct = 32'b01010100000100001101010111011110;
		#400 //-236935180.0 * -9.522148e-05 = 2488253500000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101110101011101111001111100011;
		b = 32'b10000111011011001110110010111100;
		correct = 32'b01100110101111010000100111011000;
		#400 //-7.955927e-11 * -1.7824237e-34 = 4.4635443e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100100101001001101110000000100;
		b = 32'b10100000000001011110101110110010;
		correct = 32'b01000100000111011001001000101001;
		#400 //-7.1496383e-17 * -1.1343523e-19 = 630.28375
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000001110010001001001001100011;
		b = 32'b10000010110100110010101100000001;
		correct = 32'b01111110011100110010011101111011;
		#400 //-25.071478 * -3.1028347e-37 = 8.080185e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110001111011110000000010000100;
		b = 32'b01001001000111001101100101111011;
		correct = 32'b01101000010000110000101011000101;
		#400 //2.3669613e+30 * 642455.7 = 3.6842405e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001001010001111011101000101010;
		b = 32'b00110110011111010101000111011101;
		correct = 32'b00010010010010011101011100100100;
		#400 //2.4041288e-33 * 3.7747589e-06 = 6.36896e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110001010100011001001010111101;
		b = 32'b01110011011111011111110001011000;
		correct = 32'b00111101010100110011110000111010;
		#400 //1.0377562e+30 * 2.0122822e+31 = 0.05157111
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101111000010010101011001011111;
		b = 32'b11010010010011101110110000000111;
		correct = 32'b00011100001010011110100101000111;
		#400 //-1.2490763e-10 * -222180790000.0 = 5.6218913e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010100001111001110010110110001;
		b = 32'b10110111001001110010100000111011;
		correct = 32'b01011100100100001010010110111011;
		#400 //-3245229700000.0 * -9.963343e-06 = 3.2571695e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000100011000010011101001111101;
		b = 32'b10110100001111001101010111101010;
		correct = 32'b10001111100110001010101100100001;
		#400 //2.647548e-36 * -1.7586686e-07 = -1.5054274e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011011111010000111101110001001;
		b = 32'b00100000001000100010111101001101;
		correct = 32'b01111011001101110111101100001100;
		#400 //1.3087605e+17 * 1.3737584e-19 = 9.52686e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101000001111101110010000100010;
		b = 32'b01011010111101001001011001011101;
		correct = 32'b00001100110001111100110001011100;
		#400 //1.0596587e-14 * 3.442261e+16 = 3.07838e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010010111000110011101100000100;
		b = 32'b10011101101011011111011011001111;
		correct = 32'b11110100101001110011000101001110;
		#400 //487973850000.0 * -4.6047913e-21 = -1.059709e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000010011001011100100110000000;
		b = 32'b01110000100011001000101000001011;
		correct = 32'b00010001010100010100100011110100;
		#400 //57.446777 * 3.4795828e+29 = 1.6509673e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000011101011001101011000000001;
		b = 32'b10011110001101011001100011000001;
		correct = 32'b10100100111100111010011001011011;
		#400 //1.0158384e-36 * -9.613649e-21 = -1.0566627e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101101011001111010010101101010;
		b = 32'b10110011010110001010011001010100;
		correct = 32'b01111001100010001101110000110001;
		#400 //-4.4806882e+27 * -5.0442694e-08 = 8.88273e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001011011111000101010011000011;
		b = 32'b00111000001011101001010010100101;
		correct = 32'b10010010101110010000000101101001;
		#400 //-4.8597202e-32 * 4.162327e-05 = -1.1675489e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010111110000001111111101110101;
		b = 32'b10101000111010100101000010110110;
		correct = 32'b11101110010100101101101111100000;
		#400 //424406820000000.0 * -2.6014222e-14 = -1.6314416e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000001001100010111010101110000;
		b = 32'b00011101000000110011011011000101;
		correct = 32'b10100011101011010001110010110001;
		#400 //-3.2594023e-38 * 1.736602e-21 = -1.8768849e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101111011010110111110100001011;
		b = 32'b10001100110011101000000001000011;
		correct = 32'b11100010000100011111011111001001;
		#400 //2.141755e-10 * -3.181652e-31 = -6.731582e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111011011001011110100000111101;
		b = 32'b10110100010000111000101001001111;
		correct = 32'b01000110100101100111111100011000;
		#400 //-0.0035081052 * -1.8211107e-07 = 19263.547
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111110001101101011110001010101;
		b = 32'b11111011110110001011111011100100;
		correct = 32'b01000001110101111101010010011110;
		#400 //-6.0724343e+37 * -2.2508157e+36 = 26.978817
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010110110011110000101111000111;
		b = 32'b11001010111011111000100010011011;
		correct = 32'b10001011010111010100011101110010;
		#400 //3.3450086e-25 * -7849037.5 = -4.26168e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100010010011011001000010111011;
		b = 32'b00111010000010100110100011111000;
		correct = 32'b00100111101111100001101010111110;
		#400 //2.78593e-18 * 0.0005279924 = 5.2764588e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100101100000110110010100110001;
		b = 32'b11110111100101101110011101111011;
		correct = 32'b00101101010111101110011101111101;
		#400 //-7.756208e+22 * -6.1214024e+33 = 1.267064e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010110110111011011010001011101;
		b = 32'b11011001110101100101111011100110;
		correct = 32'b00111100100001000110000100000111;
		#400 //-121883360000000.0 * -7542498400000000.0 = 0.016159547
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000100000000010010011000111111;
		b = 32'b11111101101000101110101001011011;
		correct = 32'b00000101110010101111000011101110;
		#400 //-516.5976 * -2.7068972e+37 = 1.9084492e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110001011111000010011110010110;
		b = 32'b01011100011100000001100000011101;
		correct = 32'b10010100100001100110111000000010;
		#400 //-3.6693328e-09 * 2.7032203e+17 = -1.3573933e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000100110001100110111101000000;
		b = 32'b01000111100101110010010011001000;
		correct = 32'b10111100101010000000110010101111;
		#400 //-1587.4766 * 77385.56 = -0.02051386
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000110000100101111111111111011;
		b = 32'b10011100010111100010011010011000;
		correct = 32'b11101001001010010110010111111101;
		#400 //9407.995 * -7.350352e-22 = -1.2799381e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111111111011111101101101100111;
		b = 32'b01111100100100011101011100010011;
		correct = 32'b00000010110100101000010000100001;
		#400 //1.8738831 * 6.057962e+36 = 3.0932565e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010101011001001000101001100011;
		b = 32'b11101011000110110001101001101110;
		correct = 32'b00101001101111001001101011001011;
		#400 //-15705189000000.0 * -1.8750831e+26 = 8.3757294e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100000000100010000011011001000;
		b = 32'b10101100111001110100001100110100;
		correct = 32'b10110010101000001000101000100000;
		#400 //1.2284221e-19 * -6.572876e-12 = -1.8689263e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010101010100100010101110111101;
		b = 32'b11000110110000001001111110010111;
		correct = 32'b01001110000010111010100100010011;
		#400 //-14442831000000.0 * -24655.795 = 585778370.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101001000010110011000011000100;
		b = 32'b00011111111110001000010011111100;
		correct = 32'b01001000100011110110000101010011;
		#400 //3.0906498e-14 * 1.0525209e-19 = 293642.6
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010101100111111000110000011111;
		b = 32'b10101100011100111110001001011010;
		correct = 32'b10101000101001110111100100110011;
		#400 //6.444066e-26 * -3.4658027e-12 = -1.8593286e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001110010101011101101101100000;
		b = 32'b01111001000111001011000111111111;
		correct = 32'b00010100101011101011000110011001;
		#400 //896981000.0 * 5.085053e+34 = 1.763956e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110011001111101100011001001111;
		b = 32'b11100001011010100000101001011000;
		correct = 32'b01010001010100001010110010111000;
		#400 //-1.5114724e+31 * -2.6983022e+20 = 56015684000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101000010100110011101111001011;
		b = 32'b01111011100010001110011010001000;
		correct = 32'b00101100010001011000000000010110;
		#400 //3.9900893e+24 * 1.4216562e+36 = 2.8066486e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001000110110110011100011110010;
		b = 32'b01010110010110000000000110100010;
		correct = 32'b00110010000000011110011111100000;
		#400 //448967.56 * 59375380000000.0 = 7.5615105e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001111010111000101100001100001;
		b = 32'b00110101011001110010110010110101;
		correct = 32'b00011001011101000000000111110101;
		#400 //1.08638586e-29 * 8.6119263e-07 = 1.26148996e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100101100000011110010000000110;
		b = 32'b00110011011110111011100100001100;
		correct = 32'b01110001100001000001100100000111;
		#400 //7.667395e+22 * 5.860879e-08 = 1.3082329e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110101001011110111010010110110;
		b = 32'b11111000110001000011001110010111;
		correct = 32'b00111011111001001110111001110111;
		#400 //-2.2241678e+32 * -3.1835517e+34 = 0.006986435
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010100001100101010101010000110;
		b = 32'b10111111000000011111111011000100;
		correct = 32'b10010100101011111110110010000110;
		#400 //9.020333e-27 * -0.50779366 = -1.7763776e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011100110001101101000001010010;
		b = 32'b10010100110110101100110010111110;
		correct = 32'b01000111011010001001110110110000;
		#400 //-1.315639e-21 * -2.2093131e-26 = 59549.688
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101001110111010100110111001011;
		b = 32'b10101010111011010011111010100010;
		correct = 32'b01111110011011101100110010001101;
		#400 //-3.3442497e+25 * -4.2143117e-13 = 7.935459e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011100011000001111110111011000;
		b = 32'b01000011110111110010101100111000;
		correct = 32'b00011000000000010000101110100011;
		#400 //7.444347e-22 * 446.33765 = 1.6678734e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010111100000000110010010001011;
		b = 32'b00111011100011001100001000111010;
		correct = 32'b01011011011010011000001010000110;
		#400 //282338630000000.0 * 0.0042956145 = 6.572718e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100111110011100000110100001111;
		b = 32'b01000101000101100110011111001110;
		correct = 32'b00100010001011110101101100101110;
		#400 //5.7190644e-15 * 2406.4878 = 2.3765193e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101011111110000101011111110000;
		b = 32'b01011110111110000011011000011101;
		correct = 32'b11001100100000000001000101110001;
		#400 //-6.0045775e+26 * 8.9427574e+18 = -67144584.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101010101011011000010100101111;
		b = 32'b11001101110110110110111001100011;
		correct = 32'b11011100010010100111000000011000;
		#400 //1.0488655e+26 * -460180580.0 = -2.2792477e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000011111101001000010010101100;
		b = 32'b10101101011000010100000110100111;
		correct = 32'b00010110000010101111001000000010;
		#400 //-1.4371491e-36 * -1.2804347e-11 = 1.1223915e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100110011011011001101001011001;
		b = 32'b00011111000111111001110111001000;
		correct = 32'b01000110101111101000101000001011;
		#400 //8.2435073e-16 * 3.3800073e-20 = 24389.021
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111000011101010111110010100110;
		b = 32'b10111110111010010010011100101101;
		correct = 32'b00111001000001101100010101110000;
		#400 //-5.852864e-05 * -0.455377 = 0.00012852787
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000101101101000111111000101010;
		b = 32'b00010100011110110101110111000110;
		correct = 32'b10110000101101111101000111101110;
		#400 //-1.6973464e-35 * 1.2690755e-26 = -1.3374668e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101101111100110110110000100111;
		b = 32'b10100000100111011000011010010111;
		correct = 32'b01001100110001011100101111110110;
		#400 //-2.767393e-11 * -2.6685899e-19 = 103702450.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010000101011011100110011010100;
		b = 32'b01111000101100101011110010101101;
		correct = 32'b00010111011110001110110111010100;
		#400 //23327056000.0 * 2.9001739e+34 = 8.0433303e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010011101101000110110011001000;
		b = 32'b01110011001101000011111101010101;
		correct = 32'b10100000000000000010000001000110;
		#400 //-1549838300000.0 * 1.428067e+31 = -1.08527e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001011001010000110011111110101;
		b = 32'b10100011011110110110011110001110;
		correct = 32'b11100111001010110111110000000011;
		#400 //11036661.0 * -1.3628666e-17 = -8.098123e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111101001111011111010010011100;
		b = 32'b00111011010010101110001000111001;
		correct = 32'b11000001011011111010111111101000;
		#400 //-0.046375856 * 0.0030957593 = -14.980446
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010010010010101110110001101001;
		b = 32'b11011110011110101110000101011011;
		correct = 32'b10110011010011110001000010000101;
		#400 //217887420000.0 * -4.5194576e+18 = -4.8210968e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010101111010100111011100110010;
		b = 32'b10100101100010100010110000011001;
		correct = 32'b00101111110110010011010001001000;
		#400 //-9.4699904e-26 * -2.3969066e-16 = 3.9509218e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010011010010100100101011011001;
		b = 32'b10011101111100111110001011000101;
		correct = 32'b10110100110101000101011100101110;
		#400 //2.5532887e-27 * -6.455604e-21 = -3.955151e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100001010000111100110010001101;
		b = 32'b01001011100000111101110000100111;
		correct = 32'b10010101001111100001000100111110;
		#400 //-6.633929e-19 * 17283150.0 = -3.8383796e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010011011100111100110000001111;
		b = 32'b01001001011011101001000000000010;
		correct = 32'b10001001100000101100111100000000;
		#400 //-3.077152e-27 * 977152.1 = -3.1491023e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011000010001100001101010000000;
		b = 32'b00101000010011110001001111110001;
		correct = 32'b01101111011101001110011111001010;
		#400 //871268500000000.0 * 1.1495132e-14 = 7.579456e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111100101110011111000111011011;
		b = 32'b11110100000001111111010011111110;
		correct = 32'b10001000001011110000111111101010;
		#400 //0.022698333 * -4.3086493e+31 = -5.2680854e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111010011111110010010100011011;
		b = 32'b11101001110101000111100100101110;
		correct = 32'b01010000000110011011010011100010;
		#400 //-3.3119707e+35 * -3.2108066e+25 = 10315074000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011100101111100101101110001110;
		b = 32'b00010101001100011110010011110100;
		correct = 32'b11000111000010001111011110111010;
		#400 //-1.2596812e-21 * 3.5925478e-26 = -35063.727
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100101111001111100110010011001;
		b = 32'b11111010011101110100100100101000;
		correct = 32'b10101010111011111111011110111011;
		#400 //1.368301e+23 * -3.2099528e+35 = -4.2626826e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001000100010001011101001111000;
		b = 32'b10011010011011111100001111001111;
		correct = 32'b00101101100100011111110010010100;
		#400 //-8.229041e-34 * -4.9582215e-23 = 1.6596759e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011001100111100100111111101001;
		b = 32'b11011101001010100000101000101001;
		correct = 32'b10111011111011100101100000000101;
		#400 //5570113600000000.0 * -7.657907e+17 = -0.0072736763
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001001101111000001010010100110;
		b = 32'b00100010000000001111010100111101;
		correct = 32'b00100111001110101010111011111010;
		#400 //4.527877e-33 * 1.7477063e-18 = 2.590754e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101100001011110111100011110010;
		b = 32'b00110101110100111000011001001001;
		correct = 32'b00110101110101000101111000010110;
		#400 //2.4936134e-12 * 1.5759807e-06 = 1.5822613e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000110100000001011110100100110;
		b = 32'b00011001110010001000010100101101;
		correct = 32'b00101100001001000101101110110101;
		#400 //4.842618e-35 * 2.0733305e-23 = 2.335671e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111101111010111000111000111101;
		b = 32'b01001011111100100100001000001100;
		correct = 32'b10110001011110001110101011011101;
		#400 //-0.11501739 * 31753240.0 = -3.6222254e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011100111101000100010101111100;
		b = 32'b01000000100010110000011101110101;
		correct = 32'b00011011111000001110010010111010;
		#400 //1.6164527e-21 * 4.3446603 = 3.7205503e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000111110000011100011110011110;
		b = 32'b01000010001001100110000111010010;
		correct = 32'b00000101000101010001001111001111;
		#400 //2.9156737e-34 * 41.595528 = 7.0095846e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100011101001100001100010001000;
		b = 32'b01011110001010100010011110100011;
		correct = 32'b11000100111110011110010010100111;
		#400 //-6.1278544e+21 * 3.065237e+18 = -1999.1454
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101110101000110010101100011100;
		b = 32'b00110110011110000011110010001010;
		correct = 32'b00110111101010000100010101111101;
		#400 //7.4200396e-11 * 3.6990118e-06 = 2.0059519e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110011011000000110111110000101;
		b = 32'b11001001011001111010100101010110;
		correct = 32'b01101001011110000000001111010111;
		#400 //-1.7781622e+31 * -948885.4 = 1.8739484e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101100101111011111101011110111;
		b = 32'b11001011011000100001111011110011;
		correct = 32'b01100000110101110001010101111011;
		#400 //-1.837377e+27 * -14819059.0 = 1.2398743e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011110111111100001011110101011;
		b = 32'b10110011110101001110101000110101;
		correct = 32'b10101010100110001100000101001111;
		#400 //2.6903085e-20 * -9.914621e-08 = -2.713476e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010010101011000100101001001101;
		b = 32'b01001111001101110011001101000110;
		correct = 32'b10000010111100001100000100101010;
		#400 //-1.0873043e-27 * 3073590800.0 = -3.5375701e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000110100111100101001111100000;
		b = 32'b00011011010101100100000001101111;
		correct = 32'b11101010101111010010110111000101;
		#400 //-20265.938 * 1.7722485e-22 = -1.1435156e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100011000101101001111010010;
		b = 32'b10101000100111001010001001010001;
		correct = 32'b11011011001110010101110010000110;
		#400 //907.3097 * -1.7389873e-14 = -5.21746e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000010001110110001101110101001;
		b = 32'b00010011100000001101011111011101;
		correct = 32'b01101110001110011110001000101110;
		#400 //46.77701 * 3.25246e-27 = 1.438204e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111010110110001010010010001100;
		b = 32'b01001011000110111100100111101111;
		correct = 32'b11101111001100011111111111001000;
		#400 //-5.6243676e+35 * 10209775.0 = -5.5088067e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011100010011100001000000011011;
		b = 32'b11110000000000111110110010110000;
		correct = 32'b00101011110001111110111011001111;
		#400 //-2.3200621e+17 * -1.633147e+29 = 1.4206083e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111101010111101000001100011111;
		b = 32'b11000110010110011101111100011101;
		correct = 32'b01110110100000101011100111110101;
		#400 //-1.848559e+37 * -13943.778 = 1.3257231e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000010100100100000111010000001;
		b = 32'b00000011010001110001001011111101;
		correct = 32'b00111110101110111101001001101101;
		#400 //2.1461097e-37 * 5.850264e-37 = 0.3668398
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010011101111000100101101101010;
		b = 32'b10101101110111011010000101011110;
		correct = 32'b00100101010110010111111010100010;
		#400 //-4.7532236e-27 * -2.5196453e-11 = 1.8864655e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000011011000110101011000000111;
		b = 32'b10011011111111000111011110011000;
		correct = 32'b11100110111001101000010001101000;
		#400 //227.33604 * -4.1767189e-22 = -5.4429338e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010110000101101010111101111101;
		b = 32'b10010110011001110010001110010111;
		correct = 32'b10111111001001101110010010011101;
		#400 //1.2172278e-25 * -1.8671262e-25 = -0.65192586
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110011110010100010000010111011;
		b = 32'b10011110111001101000100111100100;
		correct = 32'b11010100011000000111001110010010;
		#400 //9.4123116e-08 * -2.4409227e-20 = -3856046500000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000001010011011010011111000101;
		b = 32'b00100000100100110011000011000000;
		correct = 32'b11100000001100101101011110100101;
		#400 //-12.853459 * 2.4935029e-19 = -5.15478e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001000100011100000110000011010;
		b = 32'b00000010101100111001101001011001;
		correct = 32'b11000101010010100111100000101101;
		#400 //-8.549159e-34 * 2.6390277e-37 = -3239.511
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100000100010000100010101101000;
		b = 32'b11100001110100000110000001111110;
		correct = 32'b00111110001001110110101000111000;
		#400 //-7.855495e+19 * -4.8048447e+20 = 0.16349113
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001011010000000010111000111111;
		b = 32'b10010001110011110111001101100101;
		correct = 32'b11111000111011010010100000000001;
		#400 //12594751.0 * -3.272996e-28 = -3.8480804e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100111110101101000111000010000;
		b = 32'b11010010101101010110101100111111;
		correct = 32'b11010100100101110110000100001100;
		#400 //2.026414e+24 * -389594200000.0 = -5201346000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011010011000100110000100001000;
		b = 32'b01111011111000111000011010101000;
		correct = 32'b10011101111111101011010110100001;
		#400 //-1.5930008e+16 * 2.3627651e+36 = -6.742104e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001100111110111000101010110111;
		b = 32'b10001010111011010100010110100001;
		correct = 32'b01000001100001111011001010110111;
		#400 //-3.875616e-31 * -2.2848461e-32 = 16.962263
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000101001100001111001101011111;
		b = 32'b11010100100101101010000000101010;
		correct = 32'b10110000000101100101111011100111;
		#400 //2831.2107 * -5175457600000.0 = -5.4704546e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101000100001111011001011110010;
		b = 32'b00100001111011100101010110000101;
		correct = 32'b11000110000100011100000111100011;
		#400 //-1.5065616e-14 * 1.6150144e-18 = -9328.472
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110100101100010111010011110110;
		b = 32'b01100011010100100000010111001010;
		correct = 32'b11010000110110000100111000011011;
		#400 //-1.1247666e+32 * 3.8742334e+21 = -29031980000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100011110001100010000101110100;
		b = 32'b11001101101101011101111100010000;
		correct = 32'b01010101100010110111000101110111;
		#400 //-7.309732e+21 * -381411840.0 = 19164930000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110111010110111001100011000101;
		b = 32'b11101101010111100001011110100011;
		correct = 32'b11001001011111010001111110011000;
		#400 //4.4539514e+33 * -4.2958905e+27 = -1036793.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011011110110100110110011010010;
		b = 32'b00110101111100111000010010101010;
		correct = 32'b01100101011001011001111011100101;
		#400 //1.2296239e+17 * 1.8143521e-06 = 6.7772063e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011111111011011101110001010101;
		b = 32'b11101000011010100011000101000110;
		correct = 32'b00110111000000100000000101000000;
		#400 //-3.4279335e+19 * -4.4237708e+24 = 7.748895e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001110001100000001101101101111;
		b = 32'b11010111111110100101111101010111;
		correct = 32'b00110101101101000001000011000100;
		#400 //-738647000.0 * -550574780000000.0 = 1.3415925e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110100001000010100011000010111;
		b = 32'b10110100000110010111110111010011;
		correct = 32'b00111111100001100111110101100101;
		#400 //-1.5019792e-07 * -1.429501e-07 = 1.0507017
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000100101100010000000001101010;
		b = 32'b11101101100011101101100011011101;
		correct = 32'b00010110100111101001101011000101;
		#400 //-1416.013 * -5.5261304e+27 = 2.562395e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011001000111110010111010011000;
		b = 32'b00101100101101010100100000011100;
		correct = 32'b11101011111000001100101010100101;
		#400 //-2800359500000000.0 * 5.152335e-12 = -5.435127e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110010101110110000000001000001;
		b = 32'b10110011100000101100111110111110;
		correct = 32'b00111110101101101111101101011010;
		#400 //-2.176978e-08 * -6.091385e-08 = 0.3573864
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110100110011001100011010010110;
		b = 32'b10101111010110110010010001100010;
		correct = 32'b11000100111011110011011110100001;
		#400 //3.814245e-07 * -1.993086e-10 = -1913.7384
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100010101011100111011101100;
		b = 32'b01101111001010111001101100111110;
		correct = 32'b00010100100111110111101001100011;
		#400 //855.23315 * 5.3109613e+28 = 1.610317e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000010101100110100110111001111;
		b = 32'b10101111110011000111101001110010;
		correct = 32'b11010010011000000111101110001000;
		#400 //89.65197 * -3.7194386e-10 = -241036300000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010011110011111001010000000011;
		b = 32'b11001010110001100001101111001001;
		correct = 32'b10001000100001100001111001010001;
		#400 //5.2400097e-27 * -6491620.5 = -8.071959e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110111001111000011101011000000;
		b = 32'b00100001001111000011100111111011;
		correct = 32'b01010101100000000000000010000110;
		#400 //1.1219352e-05 * 6.3773614e-19 = 17592467000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100000011001001010000010101111;
		b = 32'b00100101010001100000001101010010;
		correct = 32'b01111010100100111100101000111111;
		#400 //6.589744e+19 * 1.7174887e-16 = 3.8368484e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100100011000011001011110101010;
		b = 32'b10110001111100100101000100111010;
		correct = 32'b11110001111011100101010010101101;
		#400 //1.6645784e+22 * -7.0523614e-09 = -2.3603136e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001100100100100000101100011010;
		b = 32'b00010101000001010110000001010011;
		correct = 32'b11110111000011000010100000010000;
		#400 //-76568780.0 * 2.6935123e-26 = -2.8427114e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010001100011110001111101101110;
		b = 32'b01001011010010110100010010010100;
		correct = 32'b01000101101101000100000001111111;
		#400 //76838450000.0 * 13321364.0 = 5768.062
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101000100100100101100110011000;
		b = 32'b01011100101101011100010101100000;
		correct = 32'b10001011010011100001110101000000;
		#400 //-1.6248111e-14 * 4.093119e+17 = -3.9696162e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101100011101101001010101100010;
		b = 32'b10001110100011101001111111011110;
		correct = 32'b01011101010111010100110010011100;
		#400 //-3.5041627e-12 * -3.515965e-30 = 9.9664324e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111010111011111101010001101001;
		b = 32'b01001110001110011011011001111101;
		correct = 32'b01101100001001010100110010100000;
		#400 //6.2263357e+35 * 778936100.0 = 7.9933845e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010011111010010101001010010111;
		b = 32'b11110111101101001010101011011101;
		correct = 32'b00011011101001010100111000101100;
		#400 //-2004226000000.0 * -7.328742e+33 = 2.7347478e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101100000010100000111100111011;
		b = 32'b00011010001110001100110111100010;
		correct = 32'b01010001001111110011111100110011;
		#400 //1.9619434e-12 * 3.821662e-23 = 51337440000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100101001111111100011101100001;
		b = 32'b01000111110010011101110101011111;
		correct = 32'b01011100111100110011010110010100;
		#400 //5.660312e+22 * 103354.74 = 5.4765863e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000001110101111101111101101111;
		b = 32'b00111001101000001000111101110110;
		correct = 32'b10000111101011000001100001110001;
		#400 //-7.929914e-38 * 0.00030624465 = -2.589405e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101100101110010110000001111000;
		b = 32'b01001000101000110101101100100001;
		correct = 32'b11100011100100010100000100111001;
		#400 //-1.7928547e+27 * 334553.03 = -5.3589554e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011111010000011100101101011011;
		b = 32'b10000101100011110101000101101111;
		correct = 32'b11011001001011010001010011001110;
		#400 //4.103755e-20 * -1.347757e-35 = -3044878000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001111101101110010100110100101;
		b = 32'b10001011101111000110010000000101;
		correct = 32'b11000011011110001110010101010000;
		#400 //1.8061234e-29 * -7.256546e-32 = -248.89575
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110001001000110101000101001000;
		b = 32'b01000101010111110010100110101010;
		correct = 32'b01101011001110110101100101001101;
		#400 //8.087091e+29 * 3570.604 = 2.2649084e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111000010010100111011110011100;
		b = 32'b11001000011000111111001001100100;
		correct = 32'b10101111011000110110001001111000;
		#400 //4.8271948e-05 * -233417.56 = -2.0680513e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010000110010011000000100000101;
		b = 32'b01000100100100000001100011000010;
		correct = 32'b11001011101100101111111010010100;
		#400 //-27045407000.0 * 1152.7737 = -23461160.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111110000111100000000110100;
		b = 32'b01011000000001010111011010010010;
		correct = 32'b10011111001110111011110011101011;
		#400 //-2.3335313e-05 * 586977200000000.0 = -3.975506e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111100001001110001100001101110;
		b = 32'b01100011011001110000000101001100;
		correct = 32'b00011000001110010010110011100000;
		#400 //0.010198696 * 4.2612913e+21 = 2.3933346e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110100101100010000110101011110;
		b = 32'b00111000100000101011011111111111;
		correct = 32'b11111011101011010101111010101101;
		#400 //-1.1222017e+32 * 6.233155e-05 = -1.8003752e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001000001000010011101010100011;
		b = 32'b10010100100011101001001110011110;
		correct = 32'b11110011000100001011111011010110;
		#400 //165098.55 * -1.439656e-26 = -1.1467916e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100000010011100100010110110011;
		b = 32'b01010010110100000001000101101011;
		correct = 32'b11001100111111011100101001100001;
		#400 //-5.945393e+19 * 446822700000.0 = -133059336.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111011001100111011100110000101;
		b = 32'b10010101011111000111011000010110;
		correct = 32'b11100101001101100011111001101110;
		#400 //0.002742381 * -5.0984148e-26 = -5.3788895e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011000011001101010100101000111;
		b = 32'b10111100111001101110001010000010;
		correct = 32'b01011010111111111100000010001011;
		#400 //-1014458860000000.0 * -0.02818418 = 3.5993911e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010000010101100010101100010001;
		b = 32'b11100010100011110001010101101010;
		correct = 32'b00101101001111111001011101001001;
		#400 //-14372586000.0 * -1.3197137e+21 = 1.0890685e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100100111110000111010000111001;
		b = 32'b10100110010000000010011010101110;
		correct = 32'b00111110001001011000000101111001;
		#400 //-1.07749744e-16 * -6.66658e-16 = 0.16162671
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111001111101000111101001010;
		b = 32'b00011000011011110100001010101101;
		correct = 32'b01101110010010111110010001011001;
		#400 //48783.29 * 3.0923689e-24 = 1.5775378e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001100010111110001110010001101;
		b = 32'b01111110111000010110011000010010;
		correct = 32'b10001100111111010110011011111101;
		#400 //-58487348.0 * 1.4980314e+38 = -3.9042806e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010001010100011000101001101000;
		b = 32'b00110101101010110001110101101100;
		correct = 32'b01011011000111001011111001101001;
		#400 //56248140000.0 * 1.2749056e-06 = 4.4119455e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110000110000111100000000101000;
		b = 32'b10110101100110000010110011000001;
		correct = 32'b10111010101001001010011100111011;
		#400 //1.4242731e-09 * -1.1337908e-06 = -0.0012562046
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010110111000001111111100011001;
		b = 32'b11110001000100010100011110001101;
		correct = 32'b00100101010001100011110001001000;
		#400 //-123693120000000.0 * -7.193892e+29 = 1.7194186e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010110110000011100101101110110;
		b = 32'b01010001001101110100001011101000;
		correct = 32'b11000101000001110101101101101101;
		#400 //-106539800000000.0 * 49193845000.0 = -2165.714
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110110100111010110110101111000;
		b = 32'b01000101101010101001011100000100;
		correct = 32'b01110000011011000011111101101000;
		#400 //1.5965057e+33 * 5458.877 = 2.9246046e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011001111110100010110010001100;
		b = 32'b10100001001001101010110001010010;
		correct = 32'b01111000010000000010000001001110;
		#400 //-8802215500000000.0 * -5.647105e-19 = 1.5587128e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010011101000010101111111111100;
		b = 32'b01010001110100010000111101110011;
		correct = 32'b00000001010001011001101110100010;
		#400 //4.073676e-27 * 112238420000.0 = 3.6294847e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011110100110111100010000110010;
		b = 32'b11001011100010001101011100100011;
		correct = 32'b10010010100100011011010000001101;
		#400 //1.6492408e-20 * -17935942.0 = -9.195172e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100000101011001011010101011001;
		b = 32'b10101001110000111110101101001011;
		correct = 32'b11110110011000011010101111100011;
		#400 //9.955961e+19 * -8.7005564e-14 = -1.1442901e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101101001110110101000111010110;
		b = 32'b01100111111111000100010010100110;
		correct = 32'b00000100101111100001011100111001;
		#400 //1.06478906e-11 * 2.3826054e+24 = 4.4690112e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110010101010110110001000110001;
		b = 32'b11101110001111001111101001110110;
		correct = 32'b01000011111010000010101001001000;
		#400 //-6.789202e+30 * -1.4621493e+28 = 464.33032
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111100011100100000110101001;
		b = 32'b00111011100000111000000100110101;
		correct = 32'b10111011100010100111011100011001;
		#400 //-1.6958295e-05 * 0.0040132054 = -0.0042256233
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011100011011101100110010010000;
		b = 32'b10000111010000001101011010001101;
		correct = 32'b11010100100111101000000111101011;
		#400 //7.9011985e-22 * -1.4507525e-34 = -5446276000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111111101111100000001110111111;
		b = 32'b01011100011000101111011110010100;
		correct = 32'b00100010110101100101001000011001;
		#400 //1.4844893 * 2.5554224e+17 = 5.809174e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011010001010001001110010111100;
		b = 32'b01110000000001010101011001000111;
		correct = 32'b00101001101000011101110100000000;
		#400 //1.1865032e+16 * 1.6506324e+29 = 7.188174e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010101110111010000110010001111;
		b = 32'b10110001001100011110100100011011;
		correct = 32'b10100100000111110000100101011010;
		#400 //8.9281003e-26 * -2.5889395e-09 = -3.448555e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011010010101100110010111001010;
		b = 32'b01101010011110000011010010111111;
		correct = 32'b00101111010111010010000101000100;
		#400 //1.5086891e+16 * 7.5015672e+25 = 2.0111651e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110000100001000000001010011100;
		b = 32'b10110101111001101011111010000010;
		correct = 32'b10111010000100100111010110001111;
		#400 //9.605006e-10 * -1.719178e-06 = -0.00055869756
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110111000001010101100110100101;
		b = 32'b11101001100001010011101011010001;
		correct = 32'b11001101000000000001110110011110;
		#400 //2.704663e+33 * -2.013311e+25 = -134339040.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110000011010011011110011001101;
		b = 32'b11110100000011011110001000011001;
		correct = 32'b10111011110100101101110111001101;
		#400 //2.8935301e+29 * -4.496458e+31 = -0.006435132
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101000001101011101001110110011;
		b = 32'b10100001011111110111100111101111;
		correct = 32'b11000110001101100011001100011110;
		#400 //1.0093423e-14 * -8.655874e-19 = -11660.779
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010010011110010011100101110011;
		b = 32'b10111111111100101000010111100110;
		correct = 32'b01010010000000111000100101110001;
		#400 //-267602670000.0 * -1.8947113 = 141236650000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100100100010110011111100011110;
		b = 32'b10111110001011101010001110000001;
		correct = 32'b11100101110011000001111010000111;
		#400 //2.0549164e+22 * -0.1705456 = -1.2049074e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010110011101100101100110110;
		b = 32'b01100100010010001010110001010110;
		correct = 32'b10010110000000111110011101110000;
		#400 //-0.0015777114 * 1.4807068e+22 = -1.0655125e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101001110110111101110110101111;
		b = 32'b01010011110110010001011001110111;
		correct = 32'b11010101100000011010001101011010;
		#400 //-3.3225203e+25 * 1864769600000.0 = -17817324000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001100101000001100101011101010;
		b = 32'b00100001001111000010101011100110;
		correct = 32'b11101010110110101100000110110110;
		#400 //-84301650.0 * 6.3753653e-19 = -1.322303e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001000100000101011100101100101;
		b = 32'b10000101101010100101011001101011;
		correct = 32'b11000010010001000111011100010011;
		#400 //7.867676e-34 * -1.6018468e-35 = -49.116283
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011111101110001111000000111011;
		b = 32'b00100111100111100101110011110101;
		correct = 32'b10110111100101010111101011100000;
		#400 //-7.832446e-20 * 4.3954594e-15 = -1.7819402e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100010111111010110001001111101;
		b = 32'b00101000100111101011001111110100;
		correct = 32'b01111001110011000101110101001111;
		#400 //2.3370615e+21 * 1.7619566e-14 = 1.3264014e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101111110111101110000100100001;
		b = 32'b10000111100101111100110111011010;
		correct = 32'b01100111101110111110111000011100;
		#400 //-4.0541528e-10 * -2.2840943e-34 = 1.7749497e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011100100001101000001001111100;
		b = 32'b11011010010100110000000001100001;
		correct = 32'b10000001101000110011001000001010;
		#400 //8.901106e-22 * -1.4847909e+16 = -5.9948546e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011011001000011110011001011000;
		b = 32'b10001011100010011000101110001011;
		correct = 32'b01001111000101101010101000100001;
		#400 //-1.3392036e-22 * -5.298044e-32 = 2527732000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000010110111100110111010110001;
		b = 32'b11011100110001101010101000000000;
		correct = 32'b10100101100011110101000001100100;
		#400 //111.216194 * -4.473517e+17 = -2.486102e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010110011110100001100001011010;
		b = 32'b01000110111010100111100110000001;
		correct = 32'b10001111000010001000011011111010;
		#400 //-2.0202523e-25 * 30012.752 = -6.731313e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010011101010100100101111011;
		b = 32'b00011101100101101100011100010011;
		correct = 32'b11011100010100000011101101101010;
		#400 //-0.0009356958 * 3.9910507e-21 = -2.3444849e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011100010111111101100110110001;
		b = 32'b10000010011010000100101110011101;
		correct = 32'b11011001011101101011000101110111;
		#400 //7.406587e-22 * -1.7066368e-37 = -4339873000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010101101010101000011011101100;
		b = 32'b00111111010111001000100001011011;
		correct = 32'b01010101110001011111001111000100;
		#400 //23437058000000.0 * 0.8614556 = 27206345000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010001010011110011000011100;
		b = 32'b01100101011000100110010100010110;
		correct = 32'b10010100010000000001110110111100;
		#400 //-0.00064811273 * 6.681997e+22 = -9.699387e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011010110001100101110100110111;
		b = 32'b10100010001101001011010010111011;
		correct = 32'b01111000000011001000001000000010;
		#400 //-2.7917268e+16 * -2.4490227e-18 = 1.139935e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000010100110111101011110100010;
		b = 32'b10010100010101111101111001110011;
		correct = 32'b10101101101110001101000001101011;
		#400 //2.289897e-37 * -1.08985964e-26 = -2.1010934e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011001011001101101000110110110;
		b = 32'b11111111001111011000111001011100;
		correct = 32'b10011001100110111101110100000111;
		#400 //4060614000000000.0 * -2.5196326e+38 = -1.6115897e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011110101000100011110010111010;
		b = 32'b00011111010011010010110010000001;
		correct = 32'b00111110110010100110110101010000;
		#400 //1.7177533e-20 * 4.344725e-20 = 0.39536524
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111000010010011101001011001;
		b = 32'b11010100011111000110000001011010;
		correct = 32'b00100010000010110011001011000000;
		#400 //-8.1794215e-06 * -4335793000000.0 = 1.886488e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101100111110010010110110001101;
		b = 32'b10010000011000000111001010100000;
		correct = 32'b01011100000011100001101001110100;
		#400 //-7.082063e-12 * -4.4264515e-29 = 1.5999413e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000011010111101111111110101110;
		b = 32'b11011110101111110001110011100101;
		correct = 32'b10100100000101010101101100011110;
		#400 //222.99875 * -6.885567e+18 = -3.2386404e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111010111001011101010111001;
		b = 32'b01101011111010110101101111101110;
		correct = 32'b10001010111100000001011001010111;
		#400 //-1.3156497e-05 * 5.690634e+26 = -2.3119563e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101010100110010110100001011111;
		b = 32'b10010101111011001011110110010110;
		correct = 32'b11010100001001011110001101000111;
		#400 //2.7250682e-13 * -9.5618755e-26 = -2849930700000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000011010010011100111011101011;
		b = 32'b10001100100011010110101001111001;
		correct = 32'b00110110001101101010100110111101;
		#400 //-5.930612e-37 * -2.178857e-31 = 2.7218914e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111110010001100000011010001;
		b = 32'b01100011011000100101001010100111;
		correct = 32'b10010011111000110001001111010011;
		#400 //-2.3931645e-05 * 4.17492e+21 = -5.7322404e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010110001001110110101100010110;
		b = 32'b11010010011011111101001010011001;
		correct = 32'b01000011001100101011011000101011;
		#400 //-46019593000000.0 * -257507600000.0 = 178.7116
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000001010011001000000010110011;
		b = 32'b00111010011010000010001110010000;
		correct = 32'b10000110011000011000010111101101;
		#400 //-3.756122e-38 * 0.0008855397 = -4.241619e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111000110001100111100111011001;
		b = 32'b11111110111101110110100100110110;
		correct = 32'b10111001010011010101110110111110;
		#400 //3.2204567e+34 * -1.644328e+38 = -0.00019585245
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000111110110010101011000111010;
		b = 32'b10110010111010010101111010001101;
		correct = 32'b00010100011011100110100110101010;
		#400 //-3.270121e-34 * -2.7167767e-08 = 1.2036768e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111011000010011001000011001100;
		b = 32'b00100010001011001010011010010001;
		correct = 32'b11011000010010111111101000101010;
		#400 //-0.0020990847 * 2.3398526e-18 = -897101200000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110110110100001110011010011111;
		b = 32'b10100101000101000000111110010111;
		correct = 32'b11010001001101001001100011000010;
		#400 //6.225731e-06 * -1.2842236e-16 = -48478560000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100100011111011010000111100011;
		b = 32'b10010100110010011110100110101101;
		correct = 32'b11001111001000001100100101110110;
		#400 //5.4997753e-17 * -2.0387982e-26 = -2697557500.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000000101011010010111000011011;
		b = 32'b00100110000100111001000110011111;
		correct = 32'b01011010000101100011011100001010;
		#400 //5.411878 * 5.1198224e-16 = 1.0570441e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111000011111111111001010000100;
		b = 32'b01110110000100001001110101000111;
		correct = 32'b01000001111000101000101011001110;
		#400 //2.0764914e+34 * 7.3328194e+32 = 28.317776
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001110011110010010000100101010;
		b = 32'b11110001111101100001111000000010;
		correct = 32'b00011100000000011001000100010000;
		#400 //-1044925060.0 * -2.4374269e+30 = 4.287001e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100101011100010101001110001011;
		b = 32'b00101110101001010111011000010010;
		correct = 32'b00110110001110101011000001011100;
		#400 //2.0931723e-16 * 7.524305e-11 = 2.7818814e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101100110110100101001010000001;
		b = 32'b01111110100011000011110010101100;
		correct = 32'b00101101110001110100010110001000;
		#400 //2.1114835e+27 * 9.320347e+37 = 2.2654559e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110110001010010001011101010111;
		b = 32'b11001001011011010100001101100111;
		correct = 32'b01101100001101100111000110111111;
		#400 //-8.573941e+32 * -971830.44 = 8.822466e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000001110010101011010010111001;
		b = 32'b01010101000101001000100110010001;
		correct = 32'b00101100001011101010110111010100;
		#400 //25.338243 * 10207410000000.0 = 2.4823381e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100000001101000010100010110100;
		b = 32'b00110001010101010010111010101110;
		correct = 32'b11101110010110000101100000001011;
		#400 //-5.1927295e+19 * 3.1022114e-09 = -1.67388e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010111111101100011011000101001;
		b = 32'b00000010100111101101011100001000;
		correct = 32'b01010100110001100110100001100010;
		#400 //1.5911049e-24 * 2.3339435e-37 = 6817238000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011100000110100001111011100;
		b = 32'b00001101111001001011101010100110;
		correct = 32'b11111101000100101110101001100001;
		#400 //-17205176.0 * 1.4096519e-30 = -1.2205266e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101000010001011010011011011000;
		b = 32'b01000111101001110011001010101011;
		correct = 32'b10100000000101110101000001110000;
		#400 //-1.0971875e-14 * 85605.336 = -1.2816812e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101110000001000110101101110011;
		b = 32'b00000110100101110110000001001010;
		correct = 32'b11100110110111111111000100011101;
		#400 //-3.010876e-11 * 5.694137e-35 = -5.2876774e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111001111011111001011000110101;
		b = 32'b01110010011010101000110000101101;
		correct = 32'b11000111000000101100000000000011;
		#400 //-1.5550069e+35 * 4.645693e+30 = -33472.01
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111101101001000011101111101101;
		b = 32'b01011010100010101101101010010110;
		correct = 32'b10100010100101110110010101110110;
		#400 //-0.080192424 * 1.9541942e+16 = -4.103606e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011101001010010010110100001100;
		b = 32'b01000100001011010110001010100011;
		correct = 32'b10011000011110011100100011110110;
		#400 //-2.2390252e-21 * 693.5412 = -3.2283955e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110101110011101010100110001100;
		b = 32'b01110001010010111101001111110101;
		correct = 32'b00000100000000011100011110101000;
		#400 //1.5397541e-06 * 1.00930716e+30 = 1.5255555e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001100101110010101111100011000;
		b = 32'b00000000111101110110001000010010;
		correct = 32'b11001011001111111101010000010000;
		#400 //-2.8560996e-31 * 2.2718549e-38 = -12571664.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000111101010011110000011100101;
		b = 32'b01000101101010011011001010100111;
		correct = 32'b11000001100000000010001011100001;
		#400 //-86977.79 * 5430.3315 = -16.01703
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100001010101100101110110101100;
		b = 32'b10001101011000001000001001111110;
		correct = 32'b11010011011101000110111011110010;
		#400 //7.2629994e-19 * -6.9182403e-31 = -1049833400000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100010110011101100010000010011;
		b = 32'b01001101000111011100100101101111;
		correct = 32'b11010101001001111011101110011100;
		#400 //-1.907079e+21 * 165451500.0 = -11526514000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000001100110111101100000000110;
		b = 32'b11001011000111010100110100000101;
		correct = 32'b10110101111111011010000011110111;
		#400 //19.48048 * -10308869.0 = -1.8896816e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000001111111111110101001101110;
		b = 32'b00101010110001000100101011011011;
		correct = 32'b00010110101001101110000100110011;
		#400 //9.4008596e-38 * 3.4868535e-13 = 2.6960867e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100011101100001001100100100110;
		b = 32'b10110000001111001110000110011110;
		correct = 32'b00110010111011110101101000100110;
		#400 //-1.9146819e-17 * -6.8714623e-10 = 2.7864257e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111110101100000000101110100010;
		b = 32'b01001010100010101011110110011100;
		correct = 32'b10110011101000100110101010110100;
		#400 //-0.34383875 * 4546254.0 = -7.563122e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110111101011111101101110000;
		b = 32'b00111100011110101011111110110100;
		correct = 32'b01000001111110110010001000101110;
		#400 //0.48043394 * 0.015304495 = 31.39169
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110000111111101101001000111110;
		b = 32'b01111001111011010110001110100000;
		correct = 32'b00110110100010010110011000111101;
		#400 //6.3090688e+29 * 1.5407437e+35 = 4.0948203e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010011111110100110110100101001;
		b = 32'b10111100111101110010100101111101;
		correct = 32'b11010110100000011011000011000111;
		#400 //2151146500000.0 * -0.03017115 = -71298130000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010000000000111101100100001101;
		b = 32'b10111100101011100000110101010010;
		correct = 32'b01010010110000011110110011010001;
		#400 //-8848160000.0 * -0.021246586 = 416450900000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101010010000110011110101010011;
		b = 32'b01100011111010010101010011100111;
		correct = 32'b00000101110101100011010100001100;
		#400 //1.7340755e-13 * 8.6084185e+21 = 2.014395e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100011101101110001100011001011;
		b = 32'b10111111000101000001111110111011;
		correct = 32'b01100100000111100011100010110110;
		#400 //-6.7550814e+21 * -0.57860917 = 1.1674688e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100000111111110000001110010000;
		b = 32'b10011111111101000010011100101101;
		correct = 32'b01000000100001011011000110100110;
		#400 //-4.3201038e-19 * -1.0340283e-19 = 4.1779356
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001101001011100001011001010011;
		b = 32'b11010000100010101000010111000010;
		correct = 32'b10111100001000001101110011110110;
		#400 //182543660.0 * -18592174000.0 = -0.009818306
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010010101100000000101101110001;
		b = 32'b00000100011001100000010111000100;
		correct = 32'b11001101110000111110110100011100;
		#400 //-1.1109982e-27 * 2.7039018e-36 = -410887040.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100111110010000101001000100100;
		b = 32'b01100001000101001011110000011001;
		correct = 32'b10000110001011000110010100000101;
		#400 //-5.560021e-15 * 1.714795e+20 = -3.2423822e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100001000000010010111100110111;
		b = 32'b10110110100111010001100001111110;
		correct = 32'b11101001110100101000010000110011;
		#400 //1.4893951e+20 * -4.681816e-06 = -3.181234e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101111000101010110001011000101;
		b = 32'b01010100010010100001010101101100;
		correct = 32'b10011010001111010011111000000100;
		#400 //-1.3586561e-10 * 3471771200000.0 = -3.913438e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110010010111101000000101000000;
		b = 32'b11100011010000111111110001110001;
		correct = 32'b01001110100100010101000111010010;
		#400 //-4.4071633e+30 * -3.6153054e+21 = 1219029200.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110101010100101001110100111100;
		b = 32'b01110111001010010100110000101001;
		correct = 32'b10111101100111110011110011110110;
		#400 //-2.6698521e+32 * 3.4337613e+33 = -0.07775299
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111001010001001011000111000011;
		b = 32'b10111100100010001001101100000111;
		correct = 32'b10111100001110000100110110110000;
		#400 //0.00018758238 * -0.016675485 = -0.011248991
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010000100011000101001111111101;
		b = 32'b11001000001001001000011101100111;
		correct = 32'b00000111110110100101100000110011;
		#400 //-5.534967e-29 * -168477.61 = 3.2852833e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011111101101010010111101010011;
		b = 32'b00000011011010100100010010011000;
		correct = 32'b11011011110001011111111000011100;
		#400 //-7.673477e-20 * 6.884516e-37 = -1.1145993e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000010101010101100100111000001;
		b = 32'b10111011001011010011101000100010;
		correct = 32'b10000110111111000110010101000110;
		#400 //2.5095056e-37 * -0.0026432355 = -9.494067e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001010101100110101001011010000;
		b = 32'b10111001111000011110010011011011;
		correct = 32'b10010000010010110011100100001100;
		#400 //1.7268224e-32 * -0.00043085855 = -4.0078638e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011010100101011111110010110000;
		b = 32'b01000010100000000010000110101000;
		correct = 32'b01010111100101011101010101001010;
		#400 //2.1108802e+16 * 64.065735 = 329486600000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111011011011100100100100100000;
		b = 32'b11111011101111001101111100011100;
		correct = 32'b10111111001000010111110100001001;
		#400 //1.2372498e+36 * -1.961354e+36 = -0.63081414
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100100010010000000110001010111;
		b = 32'b01011011111101110100001000010100;
		correct = 32'b10000111110011110001111011111000;
		#400 //-4.337854e-17 * 1.3919395e+17 = -3.11641e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100111110110001011011101101110;
		b = 32'b11011000110011101000110010101010;
		correct = 32'b01001110100001100100110011110011;
		#400 //-2.0468297e+24 * -1816828300000000.0 = 1126595000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110100000101011001111001010000;
		b = 32'b10100010110100000100110101000111;
		correct = 32'b11010000101101111110000011111110;
		#400 //1.39343e-07 * -5.6460334e-18 = -24679805000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011110100000110110011001110001;
		b = 32'b10011110111001010101101001001010;
		correct = 32'b01111111000100101010101010111000;
		#400 //-4.73419e+18 * -2.428366e-20 = 1.949537e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001000011101001100100010111011;
		b = 32'b01000010111100011011011001000010;
		correct = 32'b11000101000000011010000001111011;
		#400 //-250658.92 * 120.85597 = -2074.03
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100010001010001001111111001011;
		b = 32'b11101111101000111101010000111000;
		correct = 32'b10110010000000111011111100011011;
		#400 //7.776418e+20 * -1.0140523e+29 = -7.668656e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010000100111000101010000000010;
		b = 32'b00010010111110101011110000010010;
		correct = 32'b00111101000111111001110001101010;
		#400 //6.1660585e-29 * 1.5823581e-27 = 0.038967527
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111100111101100100110101101011;
		b = 32'b01001000000011111101011100110000;
		correct = 32'b00110100010110110010110110011010;
		#400 //0.030066213 * 147292.75 = 2.0412554e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001111101010111010000101111010;
		b = 32'b00101110010001011011100110001001;
		correct = 32'b11100000110111100011011100100010;
		#400 //-5758973000.0 * 4.4957402e-11 = -1.28098435e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111111000101011001010001111;
		b = 32'b00110011101001001000001101011010;
		correct = 32'b11000011101100000110000111111111;
		#400 //-2.7024447e-05 * 7.660738e-08 = -352.7656
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101100110000010110101101011101;
		b = 32'b11010111111010100010001110110100;
		correct = 32'b01010100010100110111101001100011;
		#400 //-1.8706375e+27 * -514878130000000.0 = 3633165600000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001000111000110010010100011101;
		b = 32'b10110101101001110010000001001100;
		correct = 32'b00010010101011011111011110111100;
		#400 //-1.3670791e-33 * -1.2451869e-06 = 1.0978906e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001111101110110001001000011111;
		b = 32'b00100110110010011110001010001000;
		correct = 32'b10101000011011010011011100001001;
		#400 //-1.8446604e-29 * 1.4008578e-15 = -1.3168077e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110110100000010010011111110100;
		b = 32'b01000100101000110010100100001000;
		correct = 32'b01110001010010101010010110100111;
		#400 //1.3097981e+33 * 1305.2822 = 1.0034597e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100011000001110100000100110110;
		b = 32'b00100000110000110001101101111111;
		correct = 32'b01000001101100010111011110101010;
		#400 //7.332174e-18 * 3.305248e-19 = 22.18343
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010011100001000111101101110101;
		b = 32'b10110010100011110011011001100010;
		correct = 32'b10100000011011001101000110111001;
		#400 //3.3443223e-27 * -1.6672121e-08 = -2.0059369e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010111001011111010100111000010;
		b = 32'b01100101100011101010011011110010;
		correct = 32'b00110001000111011001111011001111;
		#400 //193143640000000.0 * 8.4206955e+22 = 2.293678e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011100111010011110011000101100;
		b = 32'b00110110010100110010001001110000;
		correct = 32'b01100110000011011100110100001110;
		#400 //5.2669397e+17 * 3.1461495e-06 = 1.6740907e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111011011110010010011010000001;
		b = 32'b10110110110011100101111101011101;
		correct = 32'b11000100000110101000100001001111;
		#400 //0.0038017335 * -6.15038e-06 = -618.1298
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000010101000011000111010101001;
		b = 32'b11101001101101111000110101010110;
		correct = 32'b00011000011000010101001011100110;
		#400 //-80.77863 * -2.7737608e+25 = 2.9122421e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100001001011100000100001010011;
		b = 32'b11100101100110001001000010000010;
		correct = 32'b00111011000100100000001011101111;
		#400 //-2.0064583e+20 * -9.005818e+22 = 0.002227958
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001011010011111101011100100000;
		b = 32'b11001011001000011000001101101011;
		correct = 32'b10111111101001001011011011011110;
		#400 //13621024.0 * -10584939.0 = -1.2868307
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001101000011010000100000111110;
		b = 32'b00101110101111001001111101001001;
		correct = 32'b01011101101111110110100100001100;
		#400 //147882980.0 * 8.577545e-11 = 1.724071e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111100000001110100111011101111;
		b = 32'b11010001011011010011001111011011;
		correct = 32'b01101010000100100000011111110001;
		#400 //-2.810244e+36 * -63673577000.0 = 4.413517e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010111111000000000011110100000;
		b = 32'b00011010101110111111100000100101;
		correct = 32'b10111100100110001000111001001010;
		#400 //-1.4477586e-24 * 7.7742286e-23 = -0.018622536
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001111001110100010001111011010;
		b = 32'b00010011010010000110001101111001;
		correct = 32'b11111011011011011100110000011001;
		#400 //-3122911700.0 * 2.5292593e-27 = -1.23471395e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101100110101010001001101011101;
		b = 32'b11100011111000010111101000111000;
		correct = 32'b00001000011100011110101101011110;
		#400 //-6.055974e-12 * -8.3186484e+21 = 7.279997e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001111101001111001011100101100;
		b = 32'b10101000100110010100110101100011;
		correct = 32'b11100110100010111110111000010011;
		#400 //5623404500.0 * -1.7019973e-14 = -3.304003e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011111010000011001111000000111;
		b = 32'b00100001001100011100010101010110;
		correct = 32'b10111101100010110110100011101111;
		#400 //-4.1000057e-20 * 6.0231105e-19 = -0.06807124
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001100000100010111001000110110;
		b = 32'b10010101000111001110101100100111;
		correct = 32'b10110110011011010100100010011110;
		#400 //1.1204763e-31 * -3.1689452e-26 = -3.535802e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000001110100001000101101000111;
		b = 32'b11000011100011010110000100110010;
		correct = 32'b10111101101111001100111011100101;
		#400 //26.068007 * -282.75934 = -0.092191495
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110111100010000010010111011100;
		b = 32'b10111110001010100011100011111011;
		correct = 32'b11111000110011001100000100101111;
		#400 //5.5228145e+33 * -0.16623299 = -3.3223337e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111111110110101101001010101010;
		b = 32'b11000110111110110110001111011101;
		correct = 32'b10111000010111101101010111101010;
		#400 //1.709554 * -32177.932 = -5.3128148e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100101101000100011110001000110;
		b = 32'b00111111101011110100000010001001;
		correct = 32'b11100101011011001111110001100100;
		#400 //-9.57669e+22 * 1.369157 = -6.994589e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001111110110100100110100110101;
		b = 32'b00010001100011010111111000010011;
		correct = 32'b11111101110001010111110000010111;
		#400 //-7324986000.0 * 2.2323577e-28 = -3.2812778e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010101001110111010001000000100;
		b = 32'b10100011111101110011101100110010;
		correct = 32'b11110000110000100100100110101110;
		#400 //12894033000000.0 * -2.6804864e-17 = -4.8103332e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100100010111000100001101110000;
		b = 32'b01011110110000101100100100101001;
		correct = 32'b00000101000100001011111000000000;
		#400 //4.7762017e-17 * 7.0178974e+18 = 6.805745e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101101001011010000001100100010;
		b = 32'b00110000011101101010001110110100;
		correct = 32'b00111100001100111001010000010101;
		#400 //9.834607e-12 * 8.9726915e-10 = 0.0109605985
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111100110101000010010111010;
		b = 32'b11010110101000001001111101000110;
		correct = 32'b10110000011101100100010110011100;
		#400 //79113.45 * -88302970000000.0 = -8.95932e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100111100011110101001101111001;
		b = 32'b01000001110000111010110001010011;
		correct = 32'b11100101001110111000001110011100;
		#400 //-1.3536764e+24 * 24.459143 = -5.5344394e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101111100011101011000100110111;
		b = 32'b01000110100111001011011010011110;
		correct = 32'b10101000011010010001100010000011;
		#400 //-2.5955568e-10 * 20059.309 = -1.2939413e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011111011110000000010000000001;
		b = 32'b01001000111011101111101110110111;
		correct = 32'b00010110000001001101011001111000;
		#400 //5.2519355e-20 * 489437.72 = 1.073055e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011100010110111111110110110011;
		b = 32'b00110110001101100110001010010111;
		correct = 32'b00100101100110100110010001101011;
		#400 //7.278892e-22 * 2.71775e-06 = 2.6782787e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100111111101110000101100010111;
		b = 32'b01001001000011000101110101101111;
		correct = 32'b11011110011000010100011111101000;
		#400 //-2.3332582e+24 * 574934.94 = -4.0582996e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011001100011001001100111011000;
		b = 32'b01010111011111010111111111000111;
		correct = 32'b01000001100011011111110011110000;
		#400 //4946956000000000.0 * 278725240000000.0 = 17.748505
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001000011001000100110100010001;
		b = 32'b00011010111011100110111111001110;
		correct = 32'b01101100111101010001111000100010;
		#400 //233780.27 * 9.861512e-23 = 2.370633e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110011000001100110100101000001;
		b = 32'b01000000111010101110111011110100;
		correct = 32'b11110001100100100111011010111111;
		#400 //-1.0649148e+31 * 7.341669 = -1.4505077e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110110011011100001000110001011;
		b = 32'b11001011100111001100100001001101;
		correct = 32'b11101010010000100101110100001010;
		#400 //1.20715085e+33 * -20549786.0 = -5.8742743e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111111010111001101000010011000;
		b = 32'b10001111101000100001100010010010;
		correct = 32'b11101111001011100101111000011111;
		#400 //0.8625579 * -1.5983897e-29 = -5.3964177e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011011100010111100110110001001;
		b = 32'b01100001011100111110000001001101;
		correct = 32'b10111001100100101100000010111110;
		#400 //-7.870202e+16 * 2.8117009e+20 = -0.00027990894
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011000100111001000000010001110;
		b = 32'b00101100011101000011011010001110;
		correct = 32'b11101011101001000000111001000011;
		#400 //-1376607600000000.0 * 3.470477e-12 = -3.9666237e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000001000000111001100111110011;
		b = 32'b00010101111010011111100011110110;
		correct = 32'b01101010100011111111110110110110;
		#400 //8.225085 * 9.450074e-26 = 8.703725e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001101110001001010110111100001;
		b = 32'b00110011110010011001000010111001;
		correct = 32'b01011001011110011100101101011011;
		#400 //412466200.0 * 9.386117e-08 = 4394428800000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110111010001011111001110010111;
		b = 32'b10110001111100010110110011110110;
		correct = 32'b11000100110100011110011011000110;
		#400 //1.179883e-05 * -7.0264106e-09 = -1679.2117
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011100101101100010101101101011;
		b = 32'b10110100110111000010101011010111;
		correct = 32'b00100111010100111101000101101100;
		#400 //-1.2054973e-21 * -4.1009363e-07 = 2.939566e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110000010001010111101000111111;
		b = 32'b11011011011001111000111001001101;
		correct = 32'b01010100010110100101001011111110;
		#400 //-2.4446533e+29 * -6.517718e+16 = 3750781000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110011110011001000000111000010;
		b = 32'b00110101101101001111111000000010;
		correct = 32'b11111101100100001010000100111110;
		#400 //-3.2405407e+31 * 1.3484971e-06 = -2.4030756e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000000000000010101010111001011;
		b = 32'b00010101001000000101001011001101;
		correct = 32'b11101010010011101000010011001011;
		#400 //-2.0208614 * 3.237706e-26 = -6.2416454e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010111010000100110011011001111;
		b = 32'b11001001011110010111110010011000;
		correct = 32'b01001101010001110111101000010000;
		#400 //-213746820000000.0 * -1021897.5 = 209166600.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000001111001010001101000011101;
		b = 32'b10101010100110000111111010000011;
		correct = 32'b10010110110000000100110110000011;
		#400 //8.4158785e-38 * -2.708841e-13 = -3.106819e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000001010101100001110100111011;
		b = 32'b10111001001010100110011100010000;
		correct = 32'b10000111101000001101010110100010;
		#400 //3.9326564e-38 * -0.00016250857 = -2.4199686e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011110011110010110000000101110;
		b = 32'b01010001010100010100001001110000;
		correct = 32'b00001100100110001000100111001101;
		#400 //1.320184e-20 * 56172675000.0 = 2.3502244e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010101111011100001110110110011;
		b = 32'b00111000110001101111100000000100;
		correct = 32'b01011100100110010010111100011110;
		#400 //32726416000000.0 * 9.487572e-05 = 3.4493982e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110010110100010000101001110011;
		b = 32'b11010101010010111011010011000100;
		correct = 32'b10011101000000110101101000100011;
		#400 //2.4335554e-08 * -13998578000000.0 = -1.7384305e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000001100101001010000111001010;
		b = 32'b10111000001100100101101000110001;
		correct = 32'b10001000110101010101011100110010;
		#400 //5.459877e-38 * -4.2522504e-05 = -1.2839971e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001010001101101100101010010010;
		b = 32'b10101111100011111100110100010110;
		correct = 32'b01011010001000101011010010110100;
		#400 //-2994852.5 * -2.615727e-10 = 1.1449408e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011100001001100111110100100110;
		b = 32'b00100101100110001111101111000110;
		correct = 32'b11110110000010110100110011000010;
		#400 //-1.874498e+17 * 2.6538405e-16 = -7.063341e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010011011100101011011101100111;
		b = 32'b00101010000110010011001011010001;
		correct = 32'b00101000110010101100101100110100;
		#400 //3.0635119e-27 * 1.360676e-13 = 2.251463e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110010011100011100001111000001;
		b = 32'b01010110010010100001111100001111;
		correct = 32'b01011011100110010001101011111111;
		#400 //4.7886425e+30 * 55558686000000.0 = 8.619071e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001100011000101000001011010001;
		b = 32'b00011010101000010010111111111011;
		correct = 32'b11110001001100111101111110110111;
		#400 //-59378500.0 * 6.6665556e-23 = -8.9069234e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110000111111101110101011011010;
		b = 32'b11100100010001100100101110000101;
		correct = 32'b10001100001001001000110011000111;
		#400 //1.8547681e-09 * -1.4631588e+22 = -1.2676464e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111010111101000000111101001101;
		b = 32'b11110111110011000111000010110000;
		correct = 32'b01000010100110001100111001001010;
		#400 //-6.336154e+35 * -8.293079e+33 = 76.40291
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111001110001101100001000101110;
		b = 32'b01101100000101000100101110000000;
		correct = 32'b10001101001010111000111010110001;
		#400 //-0.00037910178 * 7.1711024e+26 = -5.28652e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010111110001110111001011011111;
		b = 32'b10111111100100100011110110111101;
		correct = 32'b01010111101011101001001000011111;
		#400 //-438592360000000.0 * -1.1425091 = 383885220000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100010010101001010011010010010;
		b = 32'b10011010010000111010111100000000;
		correct = 32'b01000111100010110001100100110100;
		#400 //-2.881954e-18 * -4.046642e-23 = 71218.41
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100000001011010111011101000011;
		b = 32'b10101001101011110010111100110101;
		correct = 32'b10110101111111010111110100011010;
		#400 //1.469313e-19 * -7.77975e-14 = -1.8886378e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010000111011011100011001001111;
		b = 32'b10100000011101111001000000010100;
		correct = 32'b10101111111101011110000011010101;
		#400 //9.378556e-29 * -2.0969385e-19 = -4.4724993e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100000110010100111100111100111;
		b = 32'b00001011000011010011100010111101;
		correct = 32'b11010101001101111000010100001011;
		#400 //-3.43008e-19 * 2.7198297e-32 = -12611378000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111010110001110011111101001000;
		b = 32'b10111111001111000010111010011101;
		correct = 32'b10111011000001111000011011000010;
		#400 //0.0015201354 * -0.73508626 = -0.0020679687
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010011101010001111001001100010;
		b = 32'b00100011111010111110010000111010;
		correct = 32'b00101111001101110101100100111111;
		#400 //4.264817e-27 * 2.5575409e-17 = 1.667546e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011011001011001101011001001111;
		b = 32'b10001101110111011000010011100000;
		correct = 32'b01001100110001111011110110001101;
		#400 //-1.4296753e-22 * -1.3652165e-30 = 104721510.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110001011101011111011000101011;
		b = 32'b00110111111110111000110000100111;
		correct = 32'b00111000111110100101000010110100;
		#400 //3.5792123e-09 * 2.9986795e-05 = 0.00011935961
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111101110101000001111110110001;
		b = 32'b10010111110110111100001110101001;
		correct = 32'b11100101011101110001100110000110;
		#400 //0.10357607 * -1.4201935e-24 = -7.293096e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101011011001100100011100000001;
		b = 32'b01000010001101100000000111011010;
		correct = 32'b01101000101000011111001001100110;
		#400 //2.7838824e+26 * 45.50181 = 6.11818e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010100010011100000010111011000;
		b = 32'b10101110001100100101010001101100;
		correct = 32'b01100101100100111110000010010101;
		#400 //-3539445200000.0 * -4.0547496e-11 = 8.7291335e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011100111010110100111100000110;
		b = 32'b10101101000100011010110000010011;
		correct = 32'b01101111010011101100001100100110;
		#400 //-5.2986805e+17 * -8.280504e-12 = 6.398983e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010001100111110110110010000000;
		b = 32'b00111110110111001000111000101001;
		correct = 32'b11010010001110010000101101010110;
		#400 //-85590020000.0 * 0.4307721 = -198689780000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001010110101001101001001101100;
		b = 32'b01001000011001010010000110011100;
		correct = 32'b01000001111011011100011100110111;
		#400 //6973750.0 * 234630.44 = 29.722273
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100100011011000101011011110011;
		b = 32'b10101011110101111110000101010010;
		correct = 32'b01111000000011000010000110000001;
		#400 //-1.7438788e+22 * -1.5339208e-12 = 1.1368767e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110110011000101111101011011001;
		b = 32'b00111011101100010011101101101110;
		correct = 32'b00111010001000111110110110111011;
		#400 //3.3822637e-06 * 0.005408696 = 0.0006253381
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100000010001110001000010101110;
		b = 32'b01111010111000111110001100111000;
		correct = 32'b00100100110111111001111100111101;
		#400 //5.7376625e+19 * 5.9162997e+35 = 9.6980594e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111101001010011001111101101010;
		b = 32'b01000111000111000110001100011010;
		correct = 32'b10110101100010101101010101000110;
		#400 //-0.041411795 * 40035.1 = -1.0343872e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010100010001110011100101001110;
		b = 32'b00100111101010000100011100111100;
		correct = 32'b01101100000101111000100111100010;
		#400 //3422639600000.0 * 4.67066e-15 = 7.327957e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001011010010111110101100100110;
		b = 32'b10001100010101110100100011011100;
		correct = 32'b11111110011100100111101111111111;
		#400 //13364006.0 * -1.6584923e-31 = -8.057925e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010010111010010011101001000111;
		b = 32'b10101010000110101100011010100011;
		correct = 32'b01101000010000001110000100110110;
		#400 //-500852560000.0 * -1.3746864e-13 = 3.643395e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110100001001100100011011111010;
		b = 32'b01011010110111001100011000101101;
		correct = 32'b01011000110000001100111011001101;
		#400 //5.2695365e+31 * 3.1071196e+16 = 1695955500000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100101101100111001001100111110;
		b = 32'b00011010010110110110010000000000;
		correct = 32'b11001010110100011000101001100100;
		#400 //-3.1151325e-16 * 4.5368918e-23 = -6866226.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110100000111100101000101110111;
		b = 32'b00011010110101101000010000101100;
		correct = 32'b01011000101111001110111100101000;
		#400 //1.4744533e-07 * 8.872186e-23 = 1661882800000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000011100001011111100100001100;
		b = 32'b10011001100011001111100100000001;
		correct = 32'b00101001011100110100100111100011;
		#400 //-7.874216e-37 * -1.4576233e-23 = 5.4020926e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011111111010110111010111111110;
		b = 32'b11100101100010001000110001111100;
		correct = 32'b10111001110111001011100000111011;
		#400 //3.3933493e+19 * -8.0604165e+22 = -0.00042098932
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011001010001010111111111010010;
		b = 32'b00000000001000101001111111100001;
		correct = 32'b11011001001101101000011101100111;
		#400 //-1.02104744e-23 * 3.17976e-39 = -3211082600000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000001111100011110110011111;
		b = 32'b00011001100001111011110011000000;
		correct = 32'b11010110001100110110010110000111;
		#400 //-6.9209166e-10 * 1.4034908e-23 = -49312160000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111000111001110000011100111011;
		b = 32'b01000100001100001111000010010011;
		correct = 32'b11110100001001110010000011010000;
		#400 //-3.7486476e+34 * 707.759 = -5.2965032e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100100000010011100110101101111;
		b = 32'b10100011101110100110011101101011;
		correct = 32'b00111111101111010100000010101001;
		#400 //-2.988115e-17 * -2.020996e-17 = 1.4785358
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100101000011000101010001011010;
		b = 32'b11100011111101000111101011001101;
		correct = 32'b00000000100100101111000100101011;
		#400 //-1.2171644e-16 * -9.0197086e+21 = 1.3494497e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100110100110101111000100110000;
		b = 32'b10111110111101011011011011101000;
		correct = 32'b11100111001000010110110110001111;
		#400 //3.6584678e+23 * -0.4799111 = -7.62322e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100001000001101100001111000101;
		b = 32'b10101101010011011000100010100011;
		correct = 32'b01110011001001111101101011000011;
		#400 //-1.5537315e+20 * -1.168324e-11 = 1.3298807e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101101001011010100010101010101;
		b = 32'b01000010100000110001100110011000;
		correct = 32'b10101010001010010010110001110111;
		#400 //-9.849306e-12 * 65.54999 = -1.5025642e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110100101000010011100111011;
		b = 32'b00110001100001000101101101001110;
		correct = 32'b11000100100011110100011011010001;
		#400 //-4.4153107e-06 * 3.8520858e-09 = -1146.213
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111100010010010001010001111110;
		b = 32'b01010000000110110111110000000011;
		correct = 32'b00101011101001011000100100101110;
		#400 //0.012272952 * 10434383000.0 = 1.176203e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010000110000001000100001001100;
		b = 32'b10111000001100111001100100000000;
		correct = 32'b10011000000010010011011111111010;
		#400 //7.5940645e-29 * -4.2819418e-05 = -1.7735096e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010000010101010101101110010000;
		b = 32'b00000001000100000011000110011101;
		correct = 32'b11001110101111010110010101111000;
		#400 //-4.207738e-29 * 2.648422e-38 = -1588771800.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110001000101100100011100101;
		b = 32'b01011100000000001101000101101001;
		correct = 32'b10011001101000011100000001000100;
		#400 //-2.4256817e-06 * 1.4503618e+17 = -1.6724665e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001000001001111010000100011010;
		b = 32'b10010101001011011110110011010011;
		correct = 32'b11110010011101101011101110110101;
		#400 //171652.4 * -3.5123893e-26 = -4.887055e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100100111100111101110001100100;
		b = 32'b11011011001000000001100000001100;
		correct = 32'b01001001010000101111100101101001;
		#400 //-3.5987517e+22 * -4.5062436e+16 = 798614.56
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100011100011011100101011100001;
		b = 32'b00001011100111001011111001100000;
		correct = 32'b01010111011001111001010011001000;
		#400 //1.5373173e-17 * 6.037546e-32 = 254626200000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101100001100111101000000011011;
		b = 32'b10111111001111111011101101001111;
		correct = 32'b11101100011100000001011000001001;
		#400 //8.695219e+26 * -0.74895185 = -1.160985e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010100001110010000000101110011;
		b = 32'b00010101101110001000001111011001;
		correct = 32'b00111110000000000101011100100010;
		#400 //9.340399e-27 * 7.452503e-26 = 0.12533239
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111001111011101110011001011;
		b = 32'b00110001001000010110010000111001;
		correct = 32'b01010101100101101001010010010101;
		#400 //48604.793 * 2.3485554e-09 = 20695612000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000010111010101111001101110111;
		b = 32'b00001011110011001111010110101011;
		correct = 32'b01110110100100101011101011100011;
		#400 //117.47552 * 7.894758e-32 = 1.4880192e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011001101000001001011110110111;
		b = 32'b10110111100001010110101100001010;
		correct = 32'b11100001100110100001001000101010;
		#400 //5650351000000000.0 * -1.590468e-05 = -3.5526343e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001000000001001011111001000101;
		b = 32'b00000101011100010100110011111100;
		correct = 32'b01000010000011001101010001011101;
		#400 //3.9945966e-34 * 1.1345905e-35 = 35.207386
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110110101100001010100101001000;
		b = 32'b01011010000101100100011110010011;
		correct = 32'b00011100000101100111100001110001;
		#400 //5.2649157e-06 * 1.0574986e+16 = 4.9786504e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011110101010101100001110010;
		b = 32'b01111101000111010100100000000101;
		correct = 32'b10001110001011011010000001101001;
		#400 //-27963620.0 * 1.3066421e+37 = -2.1401131e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001100101101000000000001000000;
		b = 32'b10111101010110001010011111000000;
		correct = 32'b00001110110101001011000001110011;
		#400 //-2.7733542e-31 * -0.052894354 = 5.243195e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110010011101011100011110100110;
		b = 32'b10111111010011011110111011110010;
		correct = 32'b10110010100110001100010001011010;
		#400 //1.4306272e-08 * -0.80442727 = -1.778442e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100111100010010100111111000101;
		b = 32'b11100100001100011010111010111001;
		correct = 32'b10000010110001011101010110110000;
		#400 //3.8111625e-15 * -1.3110655e+22 = -2.90692e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100000001011101100010100110101;
		b = 32'b00011010100100111000001000111111;
		correct = 32'b11000101000101111010011111110101;
		#400 //-1.4803624e-19 * 6.10082e-23 = -2426.4973
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001010010000101100011001000000;
		b = 32'b11000000110110111001111011100100;
		correct = 32'b11001000111000110000100110111110;
		#400 //3191184.0 * -6.863146 = -464973.94
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011001001010110101001111001100;
		b = 32'b10101100100110101001101000010110;
		correct = 32'b01101100000011011101100011111000;
		#400 //-3014022300000000.0 * -4.3940502e-12 = 6.859326e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000001001101111001000011110001;
		b = 32'b00101011110110110100101000011100;
		correct = 32'b00010100110101100100101111011111;
		#400 //3.3715782e-38 * 1.5581455e-12 = 2.1638404e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101010100011100010100011010011;
		b = 32'b10101111001001000010001110001011;
		correct = 32'b00111010110111011011100001000010;
		#400 //-2.5252595e-13 * -1.492834e-10 = 0.0016915875
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110001100000101110100001101101;
		b = 32'b01000111011111010111010110100010;
		correct = 32'b10101001100001000011100001010101;
		#400 //-3.8099217e-09 * 64885.633 = -5.8717496e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101111100011100111101100010110;
		b = 32'b10110011001001000000100011010010;
		correct = 32'b01111011110111100101110011000011;
		#400 //-8.819135e+28 * -3.8192248e-08 = 2.3091427e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010000011101100101000001010001;
		b = 32'b00001100101001110011110011001100;
		correct = 32'b11000011001111001000010111110101;
		#400 //-4.857682e-29 * 2.5767015e-31 = -188.52327
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101011000110001110000101101110;
		b = 32'b01110010100011000110110111001000;
		correct = 32'b10111000000010110101100110000110;
		#400 //-1.8482129e+26 * 5.562959e+30 = -3.3223558e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001110111001100100011001011101;
		b = 32'b11011011110111011100000000110101;
		correct = 32'b10110010100001001110101110011000;
		#400 //1931685500.0 * -1.2483461e+17 = -1.5473958e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001001111100000010100010110110;
		b = 32'b01000111100100010010100110111010;
		correct = 32'b11000001110100111100001110110000;
		#400 //-1967382.8 * 74323.45 = -26.47055
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001110110011100011001010001010;
		b = 32'b11101000000000101110100111110011;
		correct = 32'b10100110010010011001101110011111;
		#400 //1729709300.0 * -2.472893e+24 = -6.994679e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101101100110110000100111001110;
		b = 32'b00010101010110000100010101111111;
		correct = 32'b01010111101101111000010010111001;
		#400 //1.7625814e-11 * 4.3675675e-26 = 403561330000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100010011011011110010101100010;
		b = 32'b01000111101111111000100010010110;
		correct = 32'b00011010000111101111101111001101;
		#400 //3.2240924e-18 * 98065.17 = 3.2877037e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010001110001110101110010010001;
		b = 32'b00010011010101110000001011010110;
		correct = 32'b10111101111011010101110111111101;
		#400 //-3.1453712e-28 * 2.7138213e-27 = -0.115901925
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101010110101011011000011001011;
		b = 32'b01110110110110100111101110010110;
		correct = 32'b10110011011110100110001010001100;
		#400 //-1.2916804e+26 * 2.2156784e+33 = -5.829729e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001001100100011010010001111101;
		b = 32'b00111001101001011111000110011111;
		correct = 32'b01001111011000001010111001101111;
		#400 //1193103.6 * 0.00031651274 = 3769528000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110110111011000111110000110011;
		b = 32'b10101110010000101100000101011000;
		correct = 32'b11001000000110110110110100100110;
		#400 //7.047807e-06 * -4.4282217e-11 = -159156.6
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011111110100010010111010110101;
		b = 32'b11000100001101111100001111011001;
		correct = 32'b01011011000100011011010001001100;
		#400 //-3.0146368e+19 * -735.0601 = 4.101211e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011000100011010100111000110001;
		b = 32'b10001110000011101110001001010010;
		correct = 32'b11001001111111010010101111110000;
		#400 //3.65266e-24 * -1.761182e-30 = -2073982.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110110110011010011001001100110;
		b = 32'b01111010100001000001101000111101;
		correct = 32'b10111011110001101101001100001100;
		#400 //-2.0809435e+33 * 3.429577e+35 = -0.006067639
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000010110100010111111100111001;
		b = 32'b10011001001111111101110111101010;
		correct = 32'b10101001000010111100001011110110;
		#400 //3.0782812e-37 * -9.919284e-24 = -3.1033302e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000100000010100000001101101111;
		b = 32'b00010000111101000000000010010100;
		correct = 32'b00110010100100001100110010110100;
		#400 //1.6223399e-36 * 9.624192e-29 = 1.6856895e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010101100010010001101001111101;
		b = 32'b10011101010001001101101101101011;
		correct = 32'b11110111101100100100101101010100;
		#400 //18843357000000.0 * -2.605382e-21 = -7.232474e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011010000111011011011110000110;
		b = 32'b01000101000011100000101111111111;
		correct = 32'b01010100100011100001111011010101;
		#400 //1.1098339e+16 * 2272.7498 = 4883221000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101010100011101011100111000000;
		b = 32'b10101110111100010110010001110001;
		correct = 32'b00111011000101110101110011001101;
		#400 //-2.5353157e-13 * -1.0977253e-10 = 0.0023096085
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001111011110000110010110111011;
		b = 32'b01001001000100110100001101011000;
		correct = 32'b10000101110101111110011110111101;
		#400 //-1.22469366e-29 * 603189.5 = -2.030363e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111011000000100100010111100100;
		b = 32'b01100000101110000011000110010010;
		correct = 32'b10011001101101010000111100010010;
		#400 //-0.0019878084 * 1.061804e+20 = -1.8721048e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001000010011010010010101010100;
		b = 32'b10001011111001100100100100011111;
		correct = 32'b10111011111001000000110110010001;
		#400 //6.1733823e-34 * -8.87028e-32 = -0.006959625
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010000010100000110010000101011;
		b = 32'b00110011101100110010000101011100;
		correct = 32'b00011100000101001110100010101001;
		#400 //4.1097934e-29 * 8.341405e-08 = 4.92698e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001011111110010001011000101110;
		b = 32'b11011001100000100100010100010100;
		correct = 32'b10110001111101001011111100011100;
		#400 //32648284.0 * -4583462400000000.0 = -7.1230613e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010010100011110100110101001010;
		b = 32'b01101001110111110100110010000011;
		correct = 32'b10101000001001000100100110110000;
		#400 //-307738500000.0 * 3.3743972e+25 = -9.119807e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111111001110001010001011011111;
		b = 32'b01111001100111001001001100111010;
		correct = 32'b11000101000101101111000010011111;
		#400 //-2.4542363e+38 * 1.0162305e+35 = -2415.0388
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101000101001000100010111001011;
		b = 32'b11000000001001111010110110010100;
		correct = 32'b00100111111110101100110100000100;
		#400 //-1.8237925e-14 * -2.6199694 = 6.9611217e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010000000110000010001110011110;
		b = 32'b00001100101111100000000010010000;
		correct = 32'b01000010110011001111110000101111;
		#400 //3.0004153e-29 * 2.9274474e-31 = 102.492546
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010000000111011000001110101001;
		b = 32'b01111010101011000100011001101101;
		correct = 32'b00010100111010100001000011000110;
		#400 //10570606000.0 * 4.4725173e+35 = 2.3634578e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010110110101101010001000110101;
		b = 32'b11110100110101000110110000011011;
		correct = 32'b00100001100000010101010100011110;
		#400 //-117996080000000.0 * -1.3463862e+32 = 8.76391e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100001111101101111011110111000;
		b = 32'b10101110110110000111000110110000;
		correct = 32'b10110010100100100000110100001001;
		#400 //1.6735179e-18 * -9.842738e-11 = -1.7002565e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010100001100101101011111110001;
		b = 32'b10110011011011101111110101000011;
		correct = 32'b11100000001111111001001010111100;
		#400 //3072508300000.0 * -5.5644033e-08 = -5.521721e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101001010100010111100000100110;
		b = 32'b11001101001000000100010010000010;
		correct = 32'b01011011101001110100101110110000;
		#400 //-1.5827055e+25 * -168052770.0 = 9.417908e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111111010110011110111110110001;
		b = 32'b11110110011011000001111101110111;
		correct = 32'b01001000011011000100100001001100;
		#400 //-2.8968702e+38 * -1.1972854e+33 = 241953.19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110110000011011001110110001000;
		b = 32'b01010101110111110111001011001000;
		correct = 32'b01011111101000100011111011100101;
		#400 //7.180752e+32 * 30710510000000.0 = 2.3382067e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001000111100100111100011111101;
		b = 32'b10001010110001111011110100101000;
		correct = 32'b00111101100110110110001010100101;
		#400 //-1.4593289e-33 * -1.9234156e-32 = 0.07587174
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010101001010111011010000010111;
		b = 32'b10011000101001000100101111001100;
		correct = 32'b10111100000001011100010101011110;
		#400 //3.467524e-26 * -4.246954e-24 = -0.008164732
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001001100110000101010011010101;
		b = 32'b00010001011110010110010110100011;
		correct = 32'b11110111100111000101110101001110;
		#400 //-1247898.6 * 1.9673956e-28 = -6.3428965e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101010010100001110010001010111;
		b = 32'b11011111111001010001101010100110;
		correct = 32'b10001001111010010110101001000000;
		#400 //1.8553332e-13 * -3.301738e+19 = -5.6192627e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011110100110111100110110001100;
		b = 32'b10101000010111101110100110110000;
		correct = 32'b11110101101100101110110111001100;
		#400 //5.6133917e+18 * -1.23741485e-14 = -4.5363864e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111001000000100011111001110110;
		b = 32'b00100001100000010101110110100011;
		correct = 32'b01010111000000001101111001110011;
		#400 //0.00012421035 * 8.766165e-19 = 141692900000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100101111010110111110001001011;
		b = 32'b00010000000010101110110111110011;
		correct = 32'b01010101010110001111010111000101;
		#400 //4.0850226e-16 * 2.739901e-29 = 14909380000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000101110011111001010001011110;
		b = 32'b10111000100101111111011001110101;
		correct = 32'b10001100101011101101100011000011;
		#400 //1.9520688e-35 * -7.246147e-05 = -2.6939404e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100000011000100011110011000000;
		b = 32'b01011110100011000111000000001000;
		correct = 32'b01000001010011100011001101110011;
		#400 //6.5208463e+19 * 5.0597986e+18 = 12.887561
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110100101101000011110100110111;
		b = 32'b01101110100001110010110101110001;
		correct = 32'b00000101101010101010101101000010;
		#400 //3.3572152e-07 * 2.0917706e+28 = 1.6049633e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111010111000110000110011000110;
		b = 32'b01111000111101111010111111101111;
		correct = 32'b01000001011010101010101110000111;
		#400 //5.8945523e+35 * 4.0189553e+34 = 14.666877
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110100110010000011101000011100;
		b = 32'b01000000110111100010000111011111;
		correct = 32'b00110011011001101100000100111110;
		#400 //3.7295183e-07 * 6.9416347 = 5.37268e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110011001101101011010110100100;
		b = 32'b10111101010101110001110110011111;
		correct = 32'b00110101010110010110111101001111;
		#400 //-4.254038e-08 * -0.052518483 = 8.1000775e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110100001000010011001010100010;
		b = 32'b11111111111100001100001011000001;
		correct = 32'b11111111111100001100001011000001;
		#400 //-5.1085617e+31 * nan = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100010001010110101000010000011;
		b = 32'b00100010111000010001010100011010;
		correct = 32'b01111110110000101101100010110001;
		#400 //7.900487e+20 * 6.1008714e-18 = 1.2949768e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001001001000110011101000011111;
		b = 32'b10011011101010011011100011011101;
		correct = 32'b10101100111101100011010000000010;
		#400 //1.964774e-33 * -2.807817e-22 = -6.9975145e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100010111100100010000001011101;
		b = 32'b10111011010011010000110011101100;
		correct = 32'b10100111000101110010010011101000;
		#400 //6.5628497e-18 * -0.003128822 = -2.0975467e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101101101110000110111000001111;
		b = 32'b11100000100011000100010110010100;
		correct = 32'b10001100101010000100101110000000;
		#400 //2.0967254e-11 * -8.086118e+19 = -2.5929938e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110001101000101101111111110101;
		b = 32'b11010000001011001110111010100100;
		correct = 32'b00100000111100010001110010010010;
		#400 //-4.7402815e-09 * -11605283000.0 = 4.0845894e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100111001110111000101110000100;
		b = 32'b11011100110101110000011110101101;
		correct = 32'b11001001110111110100011100111011;
		#400 //8.8565614e+23 * -4.8420448e+17 = -1829095.4
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101011101010100000000000001101;
		b = 32'b01011110100100111101000011010100;
		correct = 32'b11001100100100110011010111100010;
		#400 //-4.1103526e+26 * 5.325623e+18 = -77180690.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110010000011001101110111001011;
		b = 32'b01111001101100110110110111101101;
		correct = 32'b00110111110010001111101011111100;
		#400 //2.790146e+30 * 1.1645634e+35 = 2.3958732e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010001001001110001000010100110;
		b = 32'b10110101111010011001111101011101;
		correct = 32'b00011010101101110001000100111100;
		#400 //-1.3179107e-28 * -1.7406234e-06 = 7.571487e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000000011000100101000000111111;
		b = 32'b11111100110001100010001000111001;
		correct = 32'b00000011000100100011010001110111;
		#400 //-3.5361478 * -8.230151e+36 = 4.296577e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011101010000001000011100101010;
		b = 32'b00111100001001100010001010101001;
		correct = 32'b01100000100101000101010110010111;
		#400 //8.6706896e+17 * 0.0101401 = 8.550892e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101111010101100101100100000100;
		b = 32'b11001101110101001001010011011011;
		correct = 32'b01100001000000010001000001000001;
		#400 //-6.6337405e+28 * -445815650.0 = 1.4880008e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100111001100011101100111000011;
		b = 32'b01110101010101000111000101011101;
		correct = 32'b10110001010101100101000010111100;
		#400 //-8.3987586e+23 * 2.6930328e+32 = -3.118699e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010111011101001110110100001010;
		b = 32'b01011101111001100100101100101001;
		correct = 32'b00111001000010000010001000000001;
		#400 //269298910000000.0 * 2.0743003e+18 = 0.00012982638
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011100001001111111000110000000;
		b = 32'b01101011010010011000101011100110;
		correct = 32'b00110000010101010101001001111010;
		#400 //1.8908741e+17 * 2.4365002e+26 = 7.7606155e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001111010100000100001010111100;
		b = 32'b11001101011000101001011111011111;
		correct = 32'b10000001011010110100100111001100;
		#400 //1.0268044e-29 * -237600240.0 = -4.321563e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101010101000011110100001011100;
		b = 32'b00101110100100100010001001000001;
		correct = 32'b10111011100011011101000100000100;
		#400 //-2.8760577e-13 * 6.645396e-11 = -0.004327895
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011000010110110110000110011101;
		b = 32'b00000001011001111000001111010011;
		correct = 32'b01010110011100101001010101000111;
		#400 //2.8354369e-24 * 4.2522578e-38 = 66680740000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011010010000010000101010110001;
		b = 32'b11010000111110011101110100101101;
		correct = 32'b01001000110001011100100001001010;
		#400 //-1.3584106e+16 * -33536174000.0 = 405058.3
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011101001101110111000111001010;
		b = 32'b11000100101100011001011010100100;
		correct = 32'b00011000000001000011100010001010;
		#400 //-2.4278676e-21 * -1420.7075 = 1.7089145e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010111111111100101111100010010;
		b = 32'b01101100011111100001000010001000;
		correct = 32'b00101011000000000010011110010010;
		#400 //559368550000000.0 * 1.2285809e+27 = 4.552965e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110101100001100000010001111000;
		b = 32'b01010010001110010011100111101110;
		correct = 32'b00100010101110010011100110000001;
		#400 //9.985079e-07 * 198885210000.0 = 5.0205235e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011110101011101100111000010001;
		b = 32'b11000110101010010101001011111000;
		correct = 32'b01010111100001000010010010101011;
		#400 //-6.298012e+18 * -21673.484 = 290586050000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011110010011011010000100110010;
		b = 32'b01110100001011001111101011000111;
		correct = 32'b00101001100110000010100011111110;
		#400 //3.7042948e+18 * 5.4819423e+31 = 6.757267e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101110011010010000000100111110;
		b = 32'b11011001010011011011111101110100;
		correct = 32'b11010100100100001111010100000111;
		#400 //1.8027877e+28 * -3619554700000000.0 = -4980689300000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100000010000111101001110010011;
		b = 32'b00010000000110110100010101101110;
		correct = 32'b01001111101000010110111010101011;
		#400 //1.6587147e-19 * 3.0621847e-29 = 5416769000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111111001101010101110011000;
		b = 32'b10101000110101011010100001000101;
		correct = 32'b11011110100010100011000100111011;
		#400 //118103.19 * -2.3720726e-14 = -4.9789026e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100011111011011000000001010011;
		b = 32'b01000001010011001000101011011000;
		correct = 32'b11100010000101001010000000010001;
		#400 //-8.76225e+21 * 12.783897 = -6.85413e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001111111110110001001000111101;
		b = 32'b01001011100101111110101001101011;
		correct = 32'b11000011110100111000101110110110;
		#400 //-8424553000.0 * 19911894.0 = -423.0915
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110010100101011001000111001010;
		b = 32'b10101011100101010011111111110101;
		correct = 32'b01000110100000000100011000101110;
		#400 //-1.741218e-08 * -1.0604838e-12 = 16419.09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011111010001010101111100001110;
		b = 32'b11100010110111110110010001001010;
		correct = 32'b10111011111000100010111001101111;
		#400 //1.4222102e+19 * -2.0604253e+21 = -0.006902508
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011101000110010000111001010010;
		b = 32'b01101110110101110100001111111010;
		correct = 32'b10101101101101100000010011000000;
		#400 //-6.893027e+17 * 3.3310728e+28 = -2.0693114e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101011010101011110101101100111;
		b = 32'b00101100000000011100010101100100;
		correct = 32'b10111110110100110000000000000100;
		#400 //-7.599949e-13 * 1.8441576e-12 = -0.4121095
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111000100011000000001011011100;
		b = 32'b10011101101110100001011001000111;
		correct = 32'b01011010010000001001110100001010;
		#400 //-6.676253e-05 * -4.9256824e-21 = 1.3553965e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011010010101011000011001100110;
		b = 32'b01001100010100011000000101001000;
		correct = 32'b11001101100000100111010011000001;
		#400 //-1.5025486e+16 * 54920480.0 = -273586200.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100000100100010111001101001111;
		b = 32'b00110110111010101001011000101101;
		correct = 32'b10101001000111101011101000110010;
		#400 //-2.464026e-19 * 6.991226e-06 = -3.5244546e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111100011001110110101100001011;
		b = 32'b11011111001010110011101001010100;
		correct = 32'b01011100101011001111111010101001;
		#400 //-4.8063667e+36 * -1.2338266e+19 = 3.8954958e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011001011111000000000110011011;
		b = 32'b10011101000110110011101000001000;
		correct = 32'b10111011110011111100110111110011;
		#400 //1.3028419e-23 * -2.054408e-21 = -0.0063416897
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100100010101110000010100010111;
		b = 32'b10110010001010100011000101101011;
		correct = 32'b00110001101000011011011010110101;
		#400 //-4.6625005e-17 * -9.906539e-09 = 4.706488e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011101100100011101111101001010;
		b = 32'b10110101101001001010101100100100;
		correct = 32'b11100111011000101100011101010000;
		#400 //1.3139002e+18 * -1.2268761e-06 = -1.0709315e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111101111101111110011011100111;
		b = 32'b11111000100011100111100011110110;
		correct = 32'b01000100110111101011100001000110;
		#400 //-4.1189779e+37 * -2.3117485e+34 = 1781.7585
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110101001101110101110110010100;
		b = 32'b00111111011011101101110001010011;
		correct = 32'b00110101010001001000010111011011;
		#400 //6.8308987e-07 * 0.9330494 = 7.3210475e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010001001010110101011101010100;
		b = 32'b01111000110000000101101000010110;
		correct = 32'b00010111111001000000100101110001;
		#400 //45994033000.0 * 3.121088e+34 = 1.4736538e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011001100010101000110101110100;
		b = 32'b10010111011000101011001111010011;
		correct = 32'b11000001100111000111010101001100;
		#400 //1.4325998e-23 * -7.325151e-25 = -19.557274
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110101011011001110100101001111;
		b = 32'b11010011010111010011011111110000;
		correct = 32'b11100001100010010001010010000001;
		#400 //3.0032083e+32 * -950126250000.0 = -3.1608518e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110110000011110001111111100100;
		b = 32'b11000110001001011101011100010111;
		correct = 32'b10101111010111001110111101010111;
		#400 //2.1327223e-06 * -10613.772 = -2.0093914e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001001101011011100010110100110;
		b = 32'b11101000101101001111001100100110;
		correct = 32'b00100000011101011101100001100010;
		#400 //-1423540.8 * -6.83609e+24 = 2.0823902e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100100000011100000000110100110;
		b = 32'b00101100011010000111011110001101;
		correct = 32'b10110111000111000110000111001001;
		#400 //-3.0792738e-17 * 3.3035547e-12 = -9.321092e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011111001001010111111111110011;
		b = 32'b10001000110111010000001110000011;
		correct = 32'b11010101101111111011001011000010;
		#400 //3.5045946e-20 * -1.3301779e-33 = -26346810000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000010011101100100110011000100;
		b = 32'b00011010001110011101001110000111;
		correct = 32'b00100111101010011010011110110111;
		#400 //1.8095256e-37 * 3.8427974e-23 = 4.708876e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100000010000000011011000010011;
		b = 32'b00111010001010000111110100100110;
		correct = 32'b10100101100100100000010110010001;
		#400 //-1.6280924e-19 * 0.000642734 = -2.5330735e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001111110100100000101110111110;
		b = 32'b10101010001001110100010011011100;
		correct = 32'b00100101001000001011101111111110;
		#400 //-2.0712122e-29 * -1.485647e-13 = 1.3941482e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101111110101100011110100000111;
		b = 32'b01111011110001010110101111101011;
		correct = 32'b00110011100010101110011101000001;
		#400 //1.3260714e+29 * 2.0501426e+36 = 6.4681906e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111000011101111010010010111110;
		b = 32'b01000101101111110110001111101110;
		correct = 32'b01110010001001011001111100011111;
		#400 //2.009123e+34 * 6124.491 = 3.280473e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111100100000100101011001111001;
		b = 32'b01100101100110111001010101110000;
		correct = 32'b00010110010101100111010110111100;
		#400 //0.015910374 * 9.184043e+22 = 1.7323933e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110100010100101101000111111;
		b = 32'b01001000110010000111010010110010;
		correct = 32'b00110101001100001011000001000011;
		#400 //0.27021977 * 410533.56 = 6.5821604e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001010100100100110101101101001;
		b = 32'b10011111000111001101001101010011;
		correct = 32'b11101010111011110000001101110110;
		#400 //4797876.5 * -3.3209088e-20 = -1.4447481e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100100100110001100001101001111;
		b = 32'b01010010010111110011000000011101;
		correct = 32'b00010001101011110011100010101111;
		#400 //6.625036e-17 * 239646230000.0 = 2.7645066e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010010001011000111000110110001;
		b = 32'b00001101010000010011011001111000;
		correct = 32'b01000100011001000111101101110110;
		#400 //5.4413766e-28 * 5.953828e-31 = 913.9291
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111011010111011101101100100011;
		b = 32'b10110011110011101100011001101011;
		correct = 32'b11000111000010010101010111100111;
		#400 //0.003385254 * -9.6287145e-08 = -35157.902
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111000010010110001001101100101;
		b = 32'b11110110001111011110010001010011;
		correct = 32'b00000001100010001110001100000111;
		#400 //-4.8417034e-05 * -9.628663e+32 = 5.028428e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010011000001110001111100110;
		b = 32'b00101110100010111111010001001110;
		correct = 32'b11001011010011011010111001011001;
		#400 //-0.00085788814 * 6.3643854e-11 = -13479513.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111000101010010101110101010111;
		b = 32'b01110010100110011010100101011001;
		correct = 32'b11000101100011010001010010100111;
		#400 //-2.748098e+34 * 6.08716e+30 = -4514.5815
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101111101001111100010001101101;
		b = 32'b01010001100100001100110010101001;
		correct = 32'b00011101100101000100110110011010;
		#400 //3.0516692e-10 * 77738615000.0 = 3.925551e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000100101100100011011000011101;
		b = 32'b10010110100010101010111011000001;
		correct = 32'b01101101101001000111101111011111;
		#400 //-1425.691 * -2.2405388e-25 = 6.3631616e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011110110111101011000010000010;
		b = 32'b00110000110101101010010110111000;
		correct = 32'b11101101100001001100101110110110;
		#400 //-8.023234e+18 * 1.5617649e-09 = -5.1372866e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101010101101100100101100100100;
		b = 32'b00110110010011110010110100010011;
		correct = 32'b00110011111000010100000011100111;
		#400 //3.2381834e-13 * 3.087164e-06 = 1.04891846e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001110011011100111010011101111;
		b = 32'b00001001001001000101010000000101;
		correct = 32'b01000100101110011011110110101011;
		#400 //2.9392066e-30 * 1.9780288e-33 = 1485.9271
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000110101001101001010110100011;
		b = 32'b10011101001110100010011101001100;
		correct = 32'b10101000111001010001011010101011;
		#400 //6.266213e-35 * -2.4637211e-21 = -2.5433938e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001101011111000010101101111111;
		b = 32'b10000100101001001001011110100010;
		correct = 32'b01001000010001000001101101110101;
		#400 //-7.770585e-31 * -3.8695467e-36 = 200813.83
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010110011010011100011010000001;
		b = 32'b10111110010111011100111111001000;
		correct = 32'b11010111100001101110011101100101;
		#400 //64259694000000.0 * -0.21661294 = -296656780000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111000101010011100111010110111;
		b = 32'b01010100000000100010100011100001;
		correct = 32'b11100100001001101111110101101101;
		#400 //-2.755284e+34 * 2236126300000.0 = -1.2321683e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111001101110010101100111001;
		b = 32'b01101010000101111110000111110110;
		correct = 32'b00011100100110100101110111011010;
		#400 //46891.223 * 4.5903717e+25 = 1.0215125e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111000000110101001011101111011;
		b = 32'b00010011111001011011110111100100;
		correct = 32'b01100011101011000100001010111110;
		#400 //3.685754e-05 * 5.7994974e-27 = 6.3552985e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111101111110000010110111111001;
		b = 32'b01011001101101111001011101000101;
		correct = 32'b00100011101011010000100000001001;
		#400 //0.121181436 * 6459530400000000.0 = 1.87601e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111000001000010100110110000000;
		b = 32'b10101000110011100100101100001110;
		correct = 32'b11001110110010000010101101000100;
		#400 //3.845757e-05 * -2.2903144e-14 = -1679139300.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110110011011010011100101100011;
		b = 32'b10111000101111000010011011000001;
		correct = 32'b11111101001000010110001001100110;
		#400 //1.2028694e+33 * -8.971757e-05 = -1.3407289e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010101111100101011011100010011;
		b = 32'b10111001101000001101101010100100;
		correct = 32'b01011011110000010010010000100010;
		#400 //-33358514000000.0 * -0.00030680478 = 1.087288e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100111100110011001110110000111;
		b = 32'b00001111101110010010101000111110;
		correct = 32'b01010111010101000110000110001000;
		#400 //4.2636822e-15 * 1.825868e-29 = 233515360000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010001010000100011010001110011;
		b = 32'b10100001110110000101010001001111;
		correct = 32'b11101110111001011101000101111111;
		#400 //52131475000.0 * -1.4659046e-18 = -3.5562666e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011101000101100101000111101011;
		b = 32'b10110001010000000001111101111100;
		correct = 32'b00101011010010000100110001100001;
		#400 //-1.9894685e-21 * -2.7957574e-09 = 7.116027e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010010111100010010111111101010;
		b = 32'b01111111011011011111010010011000;
		correct = 32'b00010011000000011011110100000111;
		#400 //517945500000.0 * 3.1629704e+38 = 1.6375287e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001101101011100000101011010111;
		b = 32'b11010101110100101001111011000000;
		correct = 32'b10110111010100111000101010001110;
		#400 //364993250.0 * -28947408000000.0 = -1.260884e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111011000111101011100100001100;
		b = 32'b00111111100010101001000110011001;
		correct = 32'b00111011000100101001110111101111;
		#400 //0.0024219183 * 1.0825683 = 0.0022371968
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010100011100011100010110111101;
		b = 32'b00110010110001010101010101101100;
		correct = 32'b01100001000111001101001100111000;
		#400 //4153618500000.0 * 2.2972664e-08 = 1.80807e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100001110111000111010000011000;
		b = 32'b11010001100000111001111101001010;
		correct = 32'b00001111110101100110001011111011;
		#400 //-1.493851e-18 * -70664140000.0 = 2.1140155e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011101000111111100001110101111;
		b = 32'b01010001111010110110101111110010;
		correct = 32'b10001010101011011011101010111111;
		#400 //-2.114464e-21 * 126391040000.0 = -1.672954e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011110101011101011000101011011;
		b = 32'b11101010010000100111101010111110;
		correct = 32'b00110011111001011111010001000010;
		#400 //-6.293971e+18 * -5.877781e+25 = 1.0708074e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011100110100001000010000111010;
		b = 32'b11000000100100011111000011011001;
		correct = 32'b01011011101101101110001000010101;
		#400 //-4.6953744e+17 * -4.5606503 = 1.0295405e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101011101110110010111010001101;
		b = 32'b01110011010100010000010110111101;
		correct = 32'b10110111111001010100000000110011;
		#400 //-4.525779e+26 * 1.6560462e+31 = -2.7328822e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100100010000001001001100111100;
		b = 32'b11100001011111011000011000101100;
		correct = 32'b01000010010000100111010010110000;
		#400 //-1.4209537e+22 * -2.922934e+20 = 48.613953
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011010011011101010101010011111;
		b = 32'b10011010011000001101100101100110;
		correct = 32'b10111111100001111101110110100011;
		#400 //4.9355073e-23 * -4.6497727e-23 = -1.0614513
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011010010001010100001011100111;
		b = 32'b11000011100001010100111101100111;
		correct = 32'b11010110001111010110011101011111;
		#400 //1.3881033e+16 * -266.62033 = -52062920000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101101111101010010001011100101;
		b = 32'b10111100110001011101010111101110;
		correct = 32'b00110000100111101001101010000101;
		#400 //-2.7868772e-11 * -0.024149861 = 1.153993e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111011000100010010001011101;
		b = 32'b10010110011000011001101011001100;
		correct = 32'b01100000100000000100111000001101;
		#400 //-1.3479116e-05 * -1.82242e-25 = 7.396273e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000111100000101001100111110000;
		b = 32'b10001001001001111101000100010111;
		correct = 32'b00111101110001110011101010010101;
		#400 //-1.9650702e-34 * -2.0200207e-33 = 0.097279705
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111011110001101001111000011100;
		b = 32'b11110101100001100111101011100000;
		correct = 32'b01000101101111010000110000010001;
		#400 //-2.0625632e+36 * -3.4094726e+32 = 6049.5083
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101001000100100011111010100000;
		b = 32'b11101110000101010000111100011010;
		correct = 32'b10111010011110110010101010100000;
		#400 //1.1049932e+25 * -1.1532881e+28 = -0.0009581242
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000011110001111100010001110010;
		b = 32'b11001110001000101010000110101000;
		correct = 32'b10110101000111010011101001011111;
		#400 //399.53473 * -682125800.0 = -5.8572e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010010010101100100111000011000;
		b = 32'b00110110000101111001011101111001;
		correct = 32'b00011011101101001111010000011001;
		#400 //6.762275e-28 * 2.2588922e-06 = 2.9936246e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000110111111101001010010011011;
		b = 32'b10011111000001000001101111010011;
		correct = 32'b01100111011101101010100110101111;
		#400 //-32586.303 * -2.7975103e-20 = 1.1648323e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100001101111000010101011011;
		b = 32'b01100010000001110111110001001000;
		correct = 32'b00100001101011010110000110101011;
		#400 //734.0837 * 6.2481646e+20 = 1.1748788e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100111100011001101100010001001;
		b = 32'b11110100100000110000111010010101;
		correct = 32'b10110010100010011000111110000000;
		#400 //1.3302514e+24 * -8.306722e+31 = -1.6014155e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100001110001000010000011010000;
		b = 32'b01000011000101111111111000000110;
		correct = 32'b01011110001001010010101101000001;
		#400 //4.5224078e+20 * 151.99228 = 2.9754195e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010111101110100110110111011000;
		b = 32'b11100100111011010101111001100110;
		correct = 32'b00110010010010010000111111100010;
		#400 //-409961880000000.0 * -3.5029444e+22 = 1.1703351e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100011100101110001011110110010;
		b = 32'b01000101111000001011110001011110;
		correct = 32'b00011101001011000001110010100010;
		#400 //1.6381488e-17 * 7191.546 = 2.2778813e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010011000011011000101010010111;
		b = 32'b00010010001101011001001000001000;
		correct = 32'b01000000010001111000111111101010;
		#400 //1.7865032e-27 * 5.7293527e-28 = 3.1181588
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110110110101010110011010110101;
		b = 32'b10001101100101001101000001000010;
		correct = 32'b11101000101101111000110111100100;
		#400 //6.3598513e-06 * -9.17134e-31 = -6.934484e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001111100101000100010110010111;
		b = 32'b10000101100001110111000010111111;
		correct = 32'b11001001100011000010000001100100;
		#400 //1.4620732e-29 * -1.2736755e-35 = -1147916.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011011100101111111001011100011;
		b = 32'b11001111000011110010111101000010;
		correct = 32'b01001100000001111101010110110010;
		#400 //-8.553956e+16 * -2402239000.0 = 35608264.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111100100110100011000111111010;
		b = 32'b01100010110101110011000010111111;
		correct = 32'b00011001001101110110111111111011;
		#400 //0.018822659 * 1.9847813e+21 = 9.4834925e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001111111011100000111101001110;
		b = 32'b11100011101011000111111010100000;
		correct = 32'b10101011101100001010011100011011;
		#400 //7987961000.0 * -6.3639285e+21 = -1.2551933e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001001101000001000100110000110;
		b = 32'b10111001110111000111011011110101;
		correct = 32'b10001111001110100110100111000111;
		#400 //3.8647925e-33 * -0.000420503 = -9.19088e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000001111010010010010001101010;
		b = 32'b10100110101101001101111011000101;
		correct = 32'b01011010101001001111111000001110;
		#400 //-29.14278 * -1.2550391e-15 = 2.3220616e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101101011001101100111011001101;
		b = 32'b01111000101111011111001001111001;
		correct = 32'b00110100000110111000100011101011;
		#400 //4.4644724e+27 * 3.0820689e+34 = 1.448531e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100000011100011001110000010110;
		b = 32'b11011100010010100011101011001011;
		correct = 32'b00000011100110001110110011100100;
		#400 //-2.0465139e-19 * -2.2769036e+17 = 8.9881445e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101000010011100100100111011010;
		b = 32'b01011100010001010101011000111001;
		correct = 32'b11001011100001011100111001110000;
		#400 //-3.8966793e+24 * 2.221815e+17 = -17538272.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001111101100010000100100010000;
		b = 32'b10111100111111100000010111000001;
		correct = 32'b11010010001100100110100111100001;
		#400 //5940322300.0 * -0.031008603 = -191570130000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111011111111010101011110001011;
		b = 32'b01101110111000000110110011101101;
		correct = 32'b00001100100100000111111000001100;
		#400 //0.007731383 * 3.4728163e+28 = 2.2262575e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011010001000101010110010001111;
		b = 32'b01100011101110011010010110001100;
		correct = 32'b10110101111000000101001001010101;
		#400 //-1.1447169e+16 * 6.849153e+21 = -1.6713262e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010011101101011101000100010000;
		b = 32'b10101101000100110000010001101100;
		correct = 32'b11100110000111100100110001000110;
		#400 //1561793100000.0 * -8.356964e-12 = -1.8688523e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100101110000010100100110101000;
		b = 32'b01010100101011001101001101010100;
		correct = 32'b10010000100011110010011110101100;
		#400 //-3.3530075e-16 * 5938239000000.0 = -5.646468e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001110010111011101100100011101;
		b = 32'b00011011011011110001010101001011;
		correct = 32'b10110010011011011000101110100001;
		#400 //-2.734489e-30 * 1.9776497e-22 = -1.3826964e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110111001010111011100010110100;
		b = 32'b01101000111100111100000101101011;
		correct = 32'b11001101101101000101100011110110;
		#400 //-3.4829257e+33 * 9.208824e+24 = -378216130.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101101000011111110011101001100;
		b = 32'b00001010101110000111101101011101;
		correct = 32'b01100001110001111011000011001010;
		#400 //8.179967e-12 * 1.776496e-32 = 4.6045513e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000100101000111011111001011111;
		b = 32'b10001101110011010000000010000110;
		correct = 32'b00110110010011000111101001010010;
		#400 //-3.8495944e-36 * -1.2634226e-30 = 3.0469569e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101101001101001101100010110000;
		b = 32'b11110000001101001101100111101100;
		correct = 32'b10111100011111111111111001000001;
		#400 //3.4980788e+27 * -2.2388301e+29 = -0.015624584
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100101100001110100111001101111;
		b = 32'b11001000010001001010111001111011;
		correct = 32'b11011100101100000001110101000010;
		#400 //7.987079e+22 * -201401.92 = -3.9657412e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111110110001011100101000000110;
		b = 32'b01110011101001010110011100101111;
		correct = 32'b11001010100110010001000000000010;
		#400 //-1.3145344e+38 * 2.620916e+31 = -5015553.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111001100000001000010000101001;
		b = 32'b10010000101110100110111011000101;
		correct = 32'b11101000001100000111100011011000;
		#400 //0.0002451253 * -7.353473e-29 = -3.3334627e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101110000111011011000011110001;
		b = 32'b01010011101011110000011011100011;
		correct = 32'b01011001111001101010010011101011;
		#400 //1.2200764e+28 * 1503469600000.0 = 8115072000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011010001100011100001000111001;
		b = 32'b10101110101000110010110010111000;
		correct = 32'b11101011000010110111000010110001;
		#400 //1.2508655e+16 * -7.4203255e-11 = -1.6857286e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111000110000111010111111000101;
		b = 32'b11001110100011100000011000111010;
		correct = 32'b10101001101100000101110100000100;
		#400 //9.331064e-05 * -1191386400.0 = -7.832106e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010010011001010001000110101111;
		b = 32'b01100000100111001110010101100000;
		correct = 32'b10110001001110101110000101111001;
		#400 //-245961050000.0 * 9.044438e+19 = -2.7194729e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011100010110111001000100111101;
		b = 32'b10001001110101111111001001000010;
		correct = 32'b01010010000000100010010101110101;
		#400 //-7.264874e-22 * -5.1987185e-33 = 139743540000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010010100101111011111000110001;
		b = 32'b00010110000000111111010000101111;
		correct = 32'b01111100000100110011001000110110;
		#400 //325865470000.0 * 1.0659146e-25 = 3.057144e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101101010001111101110110101001;
		b = 32'b10100101101000011001011000001110;
		correct = 32'b11000111000111100101001010111011;
		#400 //1.1361059e-11 * -2.803073e-16 = -40530.73
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001111101011000111110110001100;
		b = 32'b10110010010100011001111001100011;
		correct = 32'b10011100110100101010100000010010;
		#400 //1.7008868e-29 * -1.2201414e-08 = -1.3940079e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001001000111111101000000000001;
		b = 32'b11010110010011110001100010000001;
		correct = 32'b10110010010001011000110100011010;
		#400 //654592.06 * -56926038000000.0 = -1.1498992e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111001110110110011011101111110;
		b = 32'b11001000001101010001111110111100;
		correct = 32'b10110001000110101110101110001101;
		#400 //0.0004181228 * -185470.94 = -2.2543845e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111000110101010000001010010001;
		b = 32'b11100111000011110001111000111111;
		correct = 32'b10010001001111101000001001001000;
		#400 //0.000101571095 * -6.7585635e+23 = -1.5028503e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111011010010111110110010101110;
		b = 32'b11010100100111011011001011000010;
		correct = 32'b01100110001001011000010101010001;
		#400 //-1.0588367e+36 * -5418471400000.0 = 1.9541243e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000001001111111100100110010100;
		b = 32'b01010010011000010110000000010010;
		correct = 32'b10101110010110011101100100011110;
		#400 //-11.986713 * 241994860000.0 = -4.9532926e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011100010000001001011010111000;
		b = 32'b01110000101011101000100101000010;
		correct = 32'b00101011000011010011110101000000;
		#400 //2.1683565e+17 * 4.321306e+29 = 5.0178264e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001011000100010000011100001000;
		b = 32'b11000011110010110110000010100101;
		correct = 32'b00000110101101101000110101100011;
		#400 //-2.7931274e-32 * -406.75504 = 6.866854e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011110111100010110110001100100;
		b = 32'b10100011111111011111000010101111;
		correct = 32'b11111010011100110110000110110111;
		#400 //8.6981947e+18 * -2.7532248e-17 = -3.159275e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110010011010110101010101111111;
		b = 32'b00010010111101011100110110101001;
		correct = 32'b11011110111101010001100010101000;
		#400 //-1.369824e-08 * 1.5512373e-27 = -8.8305253e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100010000001100111011011010010;
		b = 32'b01000100010011011100101100010101;
		correct = 32'b00011101001001110100010011011000;
		#400 //1.822329e-18 * 823.17316 = 2.2137857e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000011010011010101100101001010;
		b = 32'b11101010111011010110011001010101;
		correct = 32'b10010111110111010111000000011000;
		#400 //205.34879 * -1.4349933e+26 = -1.4310087e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001011110010111000011111111110;
		b = 32'b00101110111001110000100000111011;
		correct = 32'b01011100011000011000011011101011;
		#400 //26677244.0 * 1.0506126e-10 = 2.5392085e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111010101100100101100100101011;
		b = 32'b01110100010111001011011111011000;
		correct = 32'b00000101110011101101101101111011;
		#400 //0.0013606896 * 6.994837e+31 = 1.9452771e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010000100001100100110110111111;
		b = 32'b00110010011000101110111111101000;
		correct = 32'b00011101100101111000000011011110;
		#400 //5.297347e-29 * 1.320948e-08 = 4.0102613e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100111101110011101010101010011;
		b = 32'b00111111100010011010010011111111;
		correct = 32'b10100111101011001100111111110001;
		#400 //-5.15791e-15 * 1.0753478 = -4.796504e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000100011111110000010111001100;
		b = 32'b00100111011001001001000011010011;
		correct = 32'b11011100100011101101000011110110;
		#400 //-1020.0906 * 3.1719866e-15 = -3.215936e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111100001011110011010101001101;
		b = 32'b10111101101001011001100100111101;
		correct = 32'b00111110000001110110110110000100;
		#400 //-0.01069386 * -0.080858685 = 0.1322537
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111010101011011111111001000;
		b = 32'b11111000001011001111101111001010;
		correct = 32'b10001110100111100010101000101001;
		#400 //54719.78 * -1.4034093e+34 = -3.8990606e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110001000101100011011100110110;
		b = 32'b11100011001111111000110000010010;
		correct = 32'b00001101010010001100001011010110;
		#400 //-2.1859257e-09 * -3.5334212e+21 = 6.1864283e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000001000001011110110111001011;
		b = 32'b00011111000001111000010101011011;
		correct = 32'b01100001011111001111111000011101;
		#400 //8.370555 * 2.869767e-20 = 2.9168064e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100110001011110011001011000010;
		b = 32'b11110010110010000010101110111101;
		correct = 32'b10110010111000000000111111111000;
		#400 //2.0683761e+23 * -7.9295844e+30 = -2.6084294e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111001011111100101100110011010;
		b = 32'b10101100111011101000000010011000;
		correct = 32'b01001100000010001000000101010011;
		#400 //-0.00024256707 * -6.7786436e-12 = 35784012.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100011101100101001111110001011;
		b = 32'b10101101000011000000101100000011;
		correct = 32'b01110110001000110100001100110011;
		#400 //-6.5900335e+21 * -7.960524e-12 = 8.278392e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100000010000110011111011000111;
		b = 32'b01001010000010110111010101111101;
		correct = 32'b00010101101100110011001111010110;
		#400 //1.6537914e-19 * 2284895.2 = 7.237931e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100110010010011111110000100011;
		b = 32'b10101111110101111101011111001101;
		correct = 32'b10110101111011111001000001001101;
		#400 //7.0077593e-16 * -3.9261608e-10 = -1.7848885e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010110000000000001101010010101;
		b = 32'b01001011010110010011100101011110;
		correct = 32'b01001010000101101111100010100001;
		#400 //35212914000000.0 * 14235998.0 = 2473512.2
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000011010111101100000100100110;
		b = 32'b10011001001111110111000101010010;
		correct = 32'b00101001100101001110111101110001;
		#400 //-6.546166e-37 * -9.8973534e-24 = 6.614057e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000000000111110011111010001011;
		b = 32'b00010011010011000110011100111101;
		correct = 32'b01101100010001110111000100010101;
		#400 //2.4881923 * 2.579932e-27 = 9.64441e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111111001000010001100100010001;
		b = 32'b11101010110111000111000010100011;
		correct = 32'b10010011101110110001010111010010;
		#400 //0.62928873 * -1.332478e+26 = -4.7226953e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111001010010010001110011110000;
		b = 32'b00110010011101100110010111000110;
		correct = 32'b11000110010100001111001101100000;
		#400 //-0.00019179634 * 1.4342225e-08 = -13372.844
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001100101101110011110110011101;
		b = 32'b00110000100110000111010010101000;
		correct = 32'b00011011100110011101100011000010;
		#400 //2.8232697e-31 * 1.1092611e-09 = 2.5451803e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001110001010110111111011011001;
		b = 32'b11110101011001011011111000011000;
		correct = 32'b00011000001111110001100010001001;
		#400 //-719304260.0 * -2.9123329e+32 = 2.4698558e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101100000001011100001011001000;
		b = 32'b11000101011001000001111100100000;
		correct = 32'b10100110000101100001101110001011;
		#400 //1.9008562e-12 * -3649.9453 = -5.207903e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101010110111110101101001000001;
		b = 32'b10110001000110001010111110010001;
		correct = 32'b10111001001110110011110111010110;
		#400 //3.9675384e-13 * -2.221871e-09 = -0.00017856745
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011010110101111001011010011000;
		b = 32'b11010001101000100100001111010001;
		correct = 32'b00001000101010100001000000110001;
		#400 //-8.9165213e-23 * -87115310000.0 = 1.0235309e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000111100000111110100111100100;
		b = 32'b00100011101011110110011001110001;
		correct = 32'b11100011010000001000011111010011;
		#400 //-67539.78 * 1.9016924e-17 = -3.551562e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101010000100110000111001010010;
		b = 32'b01101110111010110000010010011011;
		correct = 32'b10111010101000000010111101010010;
		#400 //-4.444493e+25 * 3.6367272e+28 = -0.0012221134
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101100100001010100110111100100;
		b = 32'b10111111000010001100111000010010;
		correct = 32'b01101100111110010111001100000000;
		#400 //-1.2892397e+27 * -0.5343944 = 2.4125248e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110000111011110010001110010011;
		b = 32'b10111001100001110010100101011000;
		correct = 32'b01110110111000100111011111011111;
		#400 //-5.920794e+29 * -0.0002578001 = 2.2966609e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010001100001001110000100110010;
		b = 32'b11011100011001011110110111111101;
		correct = 32'b00110100100100111111001000110100;
		#400 //-71339230000.0 * -2.5887776e+17 = 2.755711e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010100110011001100110111001101;
		b = 32'b10100001110010101100010011100110;
		correct = 32'b10110010100000010100100011010011;
		#400 //2.067991e-26 * -1.3740171e-18 = -1.5050693e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000100100011000110011101000100;
		b = 32'b10001000010011111100000001001011;
		correct = 32'b00111011101011010000001011011011;
		#400 //-3.3008676e-36 * -6.2517836e-34 = 0.0052798814
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000001010011001101100100001101;
		b = 32'b01100101110100010110011100010110;
		correct = 32'b00011010111110100110111001111110;
		#400 //12.802991 * 1.2360952e+23 = 1.03576086e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111101011011000110010001000101;
		b = 32'b10101001001100010111111010000110;
		correct = 32'b11010011101010100111100101010010;
		#400 //0.057712812 * -3.9411637e-14 = -1464359700000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111101111010100000110001101001;
		b = 32'b00000101011011000011100011010100;
		correct = 32'b01110111111111011010010011111111;
		#400 //0.11428148 * 1.1107104e-35 = 1.0289044e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110000110000000101111000011010;
		b = 32'b11101111110110110001010001000001;
		correct = 32'b01000000011000001100100101101110;
		#400 //-4.7627907e+29 * -1.35603405e+29 = 3.5122943
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011110011111010000110111000100;
		b = 32'b11111001101001101010111101010101;
		correct = 32'b00100100010000100101001011110101;
		#400 //-4.5586115e+18 * -1.0818468e+35 = 4.213731e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111001100001101011001011000001;
		b = 32'b11110000011101010001001000000010;
		correct = 32'b00001000100011001011010010011110;
		#400 //-0.00025691654 * -3.0338239e+29 = 8.468406e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011000110111111010001000110010;
		b = 32'b00011001001011111101110011000000;
		correct = 32'b00111111001000101100010100011011;
		#400 //5.7807924e-24 * 9.091868e-24 = 0.6358201
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100110011100100000111011111000;
		b = 32'b01010010110111110001100110101111;
		correct = 32'b10010011000010101110000001111101;
		#400 //-8.3980903e-16 * 479104300000.0 = -1.752873e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110001001011111001010000111010;
		b = 32'b01011011100110011011101110110100;
		correct = 32'b10010101000100100011000001100110;
		#400 //-2.5550109e-09 * 8.654411e+16 = -2.9522645e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011100000100101100111010011010;
		b = 32'b10111100011101101110100001110110;
		correct = 32'b00011111000110000011011010000100;
		#400 //-4.8574374e-22 * -0.015070071 = 3.2232346e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011110110100001000001011110001;
		b = 32'b00001000100001000001101101011110;
		correct = 32'b11010101110010100000011110000011;
		#400 //-2.2077013e-20 * 7.950895e-34 = -27766701000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001010101100010100001110110001;
		b = 32'b00001011111110110111000001001010;
		correct = 32'b01111110001101000111101011101110;
		#400 //5808600.5 * 9.6850637e-32 = 5.997483e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001101001111011111010101110110;
		b = 32'b00101011101101100110111111111000;
		correct = 32'b01100001000001010100011011110010;
		#400 //199186270.0 * 1.2962955e-12 = 1.5365807e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011101101000100001010101001000;
		b = 32'b11110010110110111010001100111100;
		correct = 32'b00101010001111001110101011000000;
		#400 //-1.459915e+18 * -8.700743e+30 = 1.67792e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111011111111000111000001100;
		b = 32'b00101100001110100100011111100111;
		correct = 32'b01011010101011111001100110111110;
		#400 //65422.047 * 2.6472104e-12 = 2.4713581e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101011011001011000000001001001;
		b = 32'b10110001101110010000000000111100;
		correct = 32'b10111001000111101100101000000111;
		#400 //8.1535175e-13 * -5.3842353e-09 = -0.00015143315
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000110001110100011110001001001;
		b = 32'b11000100110100101010100010011010;
		correct = 32'b01000000111000100101000111110101;
		#400 //-11919.071 * -1685.2688 = 7.0725045
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001001101101111010000111110101;
		b = 32'b00001011101010010001001111100010;
		correct = 32'b00111101100010110000010011010010;
		#400 //4.420795e-33 * 6.512635e-32 = 0.06788029
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011110000101101101000001100101;
		b = 32'b00110101001111010010000010111001;
		correct = 32'b10101000010011000010001110100000;
		#400 //-7.984029e-21 * 7.0455604e-07 = -1.1332e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001110011101100111000001101000;
		b = 32'b10001010100001000000011010010010;
		correct = 32'b01000011011011101110110010111110;
		#400 //-3.0375963e-30 * -1.2713609e-32 = 238.92477
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000000110010011100011010100101;
		b = 32'b11100101001111010000000110101011;
		correct = 32'b00011011000010001010010111010101;
		#400 //-6.3054986 * -5.5784877e+22 = 1.130324e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111111011000101100100100110111;
		b = 32'b11101100010101100100101111000111;
		correct = 32'b00010010100001110111010111011000;
		#400 //-0.8858828 * -1.0362719e+27 = 8.5487485e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101110010100011111001000010000;
		b = 32'b10111110100101111000010011101000;
		correct = 32'b00101111001100010101101101111001;
		#400 //-4.7736093e-11 * -0.29593587 = 1.6130554e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110001010000101010001011010011;
		b = 32'b10110100000111100010001110011000;
		correct = 32'b00111100100111011000101010001011;
		#400 //-2.832327e-09 * -1.4727846e-07 = 0.019231101
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001000000001011001001011010010;
		b = 32'b00110010000000011101000000010011;
		correct = 32'b11010101100000111011010101001101;
		#400 //-136779.28 * 7.556099e-09 = -18101838000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100011000010110110001001010101;
		b = 32'b01000111110010010001110100001000;
		correct = 32'b11011010101100010110110010000111;
		#400 //-2.571183e+21 * 102970.06 = -2.49702e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011000000111110101001000011101;
		b = 32'b00010001001110110110000110000101;
		correct = 32'b11000110010110011010101000000110;
		#400 //-2.0591725e-24 * 1.478175e-28 = -13930.506
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110011000011001111110010000101;
		b = 32'b01110001000000011111001000100111;
		correct = 32'b10000001100010101110000000001011;
		#400 //-3.2825955e-08 * 6.43461e+29 = -5.101468e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010010001010010111000010001101;
		b = 32'b00011111000000100101111111010010;
		correct = 32'b00110010101001100101101010011010;
		#400 //5.3465727e-28 * 2.760783e-20 = 1.9366144e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011110110001001111000010001111;
		b = 32'b10100001100011101101001111010101;
		correct = 32'b00111100101100000111111010011111;
		#400 //-2.08518e-20 * -9.678366e-19 = 0.021544753
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010111111111111011011010101111;
		b = 32'b01001000100010101010100100110101;
		correct = 32'b10001110111011000000110110010100;
		#400 //-1.6525105e-24 * 283977.66 = -5.8191567e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000111110111100111011001001101;
		b = 32'b01111010011101010110110100001000;
		correct = 32'b10001100111010000000101111111100;
		#400 //-113900.6 * 3.1858104e+35 = -3.5752473e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110011010001110110011101000011;
		b = 32'b01010101101010110100010001001111;
		correct = 32'b10011101000101010000011101001001;
		#400 //-4.6427214e-08 * 23538734000000.0 = -1.9723752e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111101111001100110111101111100;
		b = 32'b11010110111111111110010111111101;
		correct = 32'b01100110011001101000011011101000;
		#400 //-3.8287662e+37 * -140681630000000.0 = 2.7215822e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001110100101100010001111011011;
		b = 32'b01000101000100111101101101001011;
		correct = 32'b00001001000000011111101000001111;
		#400 //3.7012382e-30 * 2365.7058 = 1.5645387e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111111100001001010001101100;
		b = 32'b01011010101010000101101001101000;
		correct = 32'b00101100101101101110101000010100;
		#400 //123176.84 * 2.36936e+16 = 5.198739e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000111000010110000100110010000;
		b = 32'b10001111011111010001001001010011;
		correct = 32'b00110111000011001010010101101111;
		#400 //-1.0460008e-34 * -1.2477392e-29 = 8.383168e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111011001000110001010100110101;
		b = 32'b01100100011010111111000101110011;
		correct = 32'b00010110001100001111001000101111;
		#400 //0.0024884467 * 1.7409532e+22 = 1.4293586e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100010000000110110110010010001;
		b = 32'b10101101011111000101011110010001;
		correct = 32'b11110100000001010101010001000111;
		#400 //6.060866e+20 * -1.4343985e-11 = -4.2253713e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101100111000000001001100001100;
		b = 32'b01011100101001011100110000111100;
		correct = 32'b11001111101011001111110110110001;
		#400 //-2.1671146e+27 * 3.7334343e+17 = -5804614000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100001100100100100111100100001;
		b = 32'b11000011101001001000011100111011;
		correct = 32'b11011101011000111010011011010100;
		#400 //3.373658e+20 * -329.0565 = -1.025252e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111101011111100001111100110000;
		b = 32'b01101100101110110100101010110000;
		correct = 32'b01010000001011011010110001100100;
		#400 //2.1111615e+37 * 1.8113746e+27 = 11655025000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110110111111110000111001011101;
		b = 32'b10100000100111010011111101010111;
		correct = 32'b11010101110011111001110111011100;
		#400 //7.6012643e-06 * -2.663875e-19 = -28534613000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111101101111111000010010100011;
		b = 32'b11110010101100000100100011101111;
		correct = 32'b00001010100010110000111110010000;
		#400 //-0.0935147 * -6.983364e+30 = 1.3391067e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101000000111010011010001110000;
		b = 32'b10111110101010001110011010101111;
		correct = 32'b00101000111011100100010110101110;
		#400 //-8.726621e-15 * -0.32988498 = 2.6453527e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110001111010011000011111001111;
		b = 32'b11100111101000001100110100101101;
		correct = 32'b00001001101110011110010010101011;
		#400 //-6.796632e-09 * -1.5187269e+24 = 4.475217e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011011100110111100001111010111;
		b = 32'b11011011101110101011010101001001;
		correct = 32'b10111111010101011001001010111000;
		#400 //8.76879e+16 * -1.0510734e+17 = -0.83427
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110111011100101011110011000;
		b = 32'b10111010111110001000000011100001;
		correct = 32'b00111011011101011000100000111110;
		#400 //-7.10315e-06 * -0.0018959307 = 0.003746524
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000011111010011011100101011;
		b = 32'b01100001110100100111001010111010;
		correct = 32'b10001110000110100000001100100000;
		#400 //-9.211926e-10 * 4.852604e+20 = -1.898347e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010010110110101110101011010000;
		b = 32'b00101111100111110010011101110100;
		correct = 32'b10100010101100000001000010001010;
		#400 //-1.381562e-27 * 2.8949965e-10 = -4.7722407e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110110100011011100101000110011;
		b = 32'b11100010111111100011100011111101;
		correct = 32'b11010011000011101100011111111010;
		#400 //1.4379198e+33 * -2.3447897e+21 = -613240400000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001111110001101111101100010010;
		b = 32'b10000111111110100010011100001000;
		correct = 32'b01000111010010111010000111010001;
		#400 //-1.9621016e-29 * -3.763876e-34 = 52129.816
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110010011100011100100100000001;
		b = 32'b11111111001110000010111011110110;
		correct = 32'b00110010101010000000011111100110;
		#400 //-4.7890487e+30 * -2.4482179e+38 = 1.9561366e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011111100110001110111001010100;
		b = 32'b11010010100100111010000000101001;
		correct = 32'b11001100100001001001100110011100;
		#400 //2.2039675e+19 * -317023620000.0 = -69520610.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001100101111010011110111101000;
		b = 32'b00000111101110010010101111001110;
		correct = 32'b11000100100000101101000001011011;
		#400 //-2.915732e-31 * 2.7861452e-34 = -1046.5111
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101001000101101101101001110100;
		b = 32'b01010111100010000001111101010111;
		correct = 32'b11010001000011011101101000010111;
		#400 //-1.1398156e+25 * 299336370000000.0 = -38078083000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001000010000011000011111000000;
		b = 32'b00001111111101100110100011110100;
		correct = 32'b10110111110010010000111111110001;
		#400 //-5.82384e-34 * 2.42979e-29 = -2.396849e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100101100011100000001001110010;
		b = 32'b00110110010011000001001111110100;
		correct = 32'b01101110101100100010001111010111;
		#400 //8.382764e+22 * 3.0409983e-06 = 2.756583e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011000101111010101000101010011;
		b = 32'b00001100001011111001101101101111;
		correct = 32'b01001100000010011111111001011100;
		#400 //4.893747e-24 * 1.3528284e-31 = 36174190.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110010001100001111110110101010;
		b = 32'b01000111010010010001010110100101;
		correct = 32'b00101010011000010101001110010001;
		#400 //1.0302225e-08 * 51477.645 = 2.0013007e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110001000001010101110011001011;
		b = 32'b01100100010111011000000011100110;
		correct = 32'b11001100000110100010000111001111;
		#400 //-6.60379e+29 * 1.6344074e+22 = -40404796.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111001001010000100100011001101;
		b = 32'b10100010110111110100110000000100;
		correct = 32'b11010101110000001110111000111001;
		#400 //0.00016048849 * -6.0524756e-18 = -26516174000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110001110001011010011100110100;
		b = 32'b11001011101100111101111110111001;
		correct = 32'b00100101100011001010011011100001;
		#400 //-5.7524634e-09 * -23576434.0 = 2.439921e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111110111010100011111000101;
		b = 32'b00101111100111101110000011110101;
		correct = 32'b11000111101100100100011000001011;
		#400 //-2.6378673e-05 * 2.8899874e-10 = -91276.086
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101011100011001011010001101001;
		b = 32'b11010101011000111100110001011100;
		correct = 32'b01010101100111100001111111001001;
		#400 //-3.4020316e+26 * -15654179000000.0 = 21732420000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101000101111111001111010110001;
		b = 32'b10010011100100110000010101011000;
		correct = 32'b01010100101001101101010000111001;
		#400 //-2.1274081e-14 * -3.7113286e-27 = 5732200600000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100100001110001100000110100100;
		b = 32'b11000110100100110010111111001010;
		correct = 32'b00011101001000001010110000011011;
		#400 //-4.006266e-17 * -18839.895 = 2.12648e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001010100010111011001100101001;
		b = 32'b00111101011110110000111010000100;
		correct = 32'b10001100100011100111001101010110;
		#400 //-1.3452606e-32 * 0.06129314 = -2.194798e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001111011111001001001110100111;
		b = 32'b00000110110010001100010001100001;
		correct = 32'b11001000001000010000100000010000;
		#400 //-1.2452996e-29 * 7.552019e-35 = -164896.25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010101000111010101001011101011;
		b = 32'b00110000011001100101010001010101;
		correct = 32'b10100100001011101101101110011111;
		#400 //-3.1771308e-26 * 8.3793356e-10 = -3.7916262e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111011001100000101010000111110;
		b = 32'b11110001110000100011101001010110;
		correct = 32'b00001000111010000110100010011111;
		#400 //-0.002690568 * -1.9235397e+30 = 1.3987588e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010101001011001011011000111000;
		b = 32'b00001110000101001100010000111000;
		correct = 32'b01000110100101001001101001001110;
		#400 //3.487887e-26 * 1.8336884e-30 = 19021.152
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111101010101001111100100001101;
		b = 32'b10011100101110011010001100100010;
		correct = 32'b11100000000100101101100100101111;
		#400 //0.051995326 * -1.2284442e-21 = -4.232616e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101011101011110101001001001010;
		b = 32'b00010000000101110001100100011010;
		correct = 32'b11011011000101001000010100111001;
		#400 //-1.2457338e-12 * 2.9798837e-29 = -4.1804776e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011101111000100110011001010010;
		b = 32'b11110010010010111000000011001000;
		correct = 32'b00101011000011100110011011001111;
		#400 //-2.0392271e+18 * -4.0307932e+30 = 5.059121e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011000000110001111001011001;
		b = 32'b01001011000011010001110001010111;
		correct = 32'b10111111011011011101111101011000;
		#400 //-8592985.0 * 9247831.0 = -0.9291892
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000110000100010100001011110011;
		b = 32'b10000001110001111101110011011001;
		correct = 32'b01000011101110100000111111111111;
		#400 //-2.7320655e-35 * -7.3417956e-38 = 372.12497
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010011000000000111100100100110;
		b = 32'b00010100100110100100111000101100;
		correct = 32'b11111101110101010010010010101101;
		#400 //-551788350000.0 * 1.558086e-26 = -3.54145e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010011111011010101000000010101;
		b = 32'b10100110100111011001000101110101;
		correct = 32'b10101100110000001100011111000001;
		#400 //5.9906178e-27 * -1.093349e-15 = -5.4791453e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100111001011100111111110101000;
		b = 32'b11001101001001001100111010111110;
		correct = 32'b00011001100001111000011011010110;
		#400 //-2.4216553e-15 * -172813280.0 = 1.4013133e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100110011110110111011001010110;
		b = 32'b10000111111110001101100011100111;
		correct = 32'b11011110000000010101100001010110;
		#400 //8.7243494e-16 * -3.7442376e-34 = -2.3300735e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000110010000110011001010001111;
		b = 32'b01010001100100010011010111011010;
		correct = 32'b00110100001011000001000000001010;
		#400 //12492.64 * 77959220000.0 = 1.6024583e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000000111010111110001011011100;
		b = 32'b00010100101111001101010010011101;
		correct = 32'b10101011100111111110010110100000;
		#400 //-2.1662723e-38 * 1.906701e-26 = -1.1361363e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001011110001100000110110101001;
		b = 32'b01001010000010011001001110010110;
		correct = 32'b10000001001110000100010001100100;
		#400 //-7.628738e-32 * 2254053.5 = -3.384453e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101010110110001000001000001011;
		b = 32'b11100101010100010101110110101000;
		correct = 32'b01000101000001000101110111010010;
		#400 //-1.3087104e+26 * -6.179389e+22 = 2117.8638
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100111111111011000110111000101;
		b = 32'b00100100011000101100001100100110;
		correct = 32'b11000011000011110001111101111000;
		#400 //-7.0375313e-15 * 4.9171235e-17 = -143.12292
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111111111010111101011011011001;
		b = 32'b01000101110000000001001001001111;
		correct = 32'b01111111111010111101011011011001;
		#400 //nan * 6146.2886 = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101010111011011101101101011100;
		b = 32'b00101011000000010110001111001110;
		correct = 32'b11111111011010110100110101001001;
		#400 //-1.4377566e+26 * 4.5968513e-13 = -3.1276987e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011101011000110101000100110001;
		b = 32'b00000001101011000101010100101010;
		correct = 32'b11011011001010001101011011110110;
		#400 //-3.0085175e-21 * 6.3305026e-38 = -4.752415e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011010000011101101110001000011;
		b = 32'b10010111010011110011010100011011;
		correct = 32'b11000010001100001000000000101111;
		#400 //2.9542838e-23 * -6.6952336e-25 = -44.12518
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111000000100000100000011001;
		b = 32'b10001010100111000010100011100011;
		correct = 32'b01101011110101010010101011000000;
		#400 //-7.750489e-06 * -1.5037633e-32 = 5.1540616e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010001001100011100100000001100;
		b = 32'b10001001111110100001101001010011;
		correct = 32'b01000110101101011111100100101101;
		#400 //-1.4024482e-28 * -6.0210066e-33 = 23292.588
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111110000010100100111000011101;
		b = 32'b11110111000000111011110101101111;
		correct = 32'b00000110100001100110000011110111;
		#400 //-0.1350636 * -2.672004e+33 = 5.0547675e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111000110100011000001110111001;
		b = 32'b11011000100111101101101100010110;
		correct = 32'b01011111101010001101000110100011;
		#400 //-3.3995678e+34 * -1397310400000000.0 = 2.4329367e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100100110011000110001001000011;
		b = 32'b01000101001100000000010111011011;
		correct = 32'b01011111000101001001111110011100;
		#400 //3.016173e+22 * 2816.366 = 1.070945e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111100100101110100110100010100;
		b = 32'b01101101100110000100110100100001;
		correct = 32'b11001110011111100101000110011100;
		#400 //-6.284801e+36 * 5.8918706e+27 = -1066690300.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111101100111110000110110101010;
		b = 32'b01110100101001101000010100111001;
		correct = 32'b11001000011101001000010101000100;
		#400 //-2.6427275e+37 * 1.0554484e+32 = -250389.06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110100011110110000101000110010;
		b = 32'b11100100011110010001100111001101;
		correct = 32'b00001111100000001111111100010010;
		#400 //-2.3379906e-07 * -1.8380394e+22 = 1.2720024e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010011000110101010111011101110;
		b = 32'b01001001011100000001101101100010;
		correct = 32'b11001001001001001110110000001011;
		#400 //-664359800000.0 * 983478.1 = -675520.7
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011011100101101101101010011010;
		b = 32'b00111010000000100001000001000000;
		correct = 32'b00100001000101000111010111101001;
		#400 //2.4956686e-22 * 0.0004961528 = 5.0300403e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101000011101100010100101110010;
		b = 32'b11100000000011111101101111011011;
		correct = 32'b00000111110110110000011001111100;
		#400 //-1.366473e-14 * -4.146448e+19 = 3.2955269e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100001010000110010101011000000;
		b = 32'b10100000111111011011101010110101;
		correct = 32'b10111111110001001110100111100000;
		#400 //6.612515e-19 * -4.298342e-19 = -1.5383873
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111100001111001110101111001111;
		b = 32'b01001010000010011110001111010001;
		correct = 32'b01110001101011110101111100000000;
		#400 //3.9237383e+36 * 2259188.2 = 1.7367912e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001110101010100111111011110100;
		b = 32'b00011011111101110100111010001101;
		correct = 32'b01110010001100000111110100110011;
		#400 //1430223400.0 * 4.0913485e-22 = 3.495726e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011000111101010000101111111100;
		b = 32'b10011110111011101000011110100100;
		correct = 32'b01111001100000110111111101000100;
		#400 //-2155454600000000.0 * -2.525533e-20 = 8.534652e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001011011000111010101110111101;
		b = 32'b10001011001101000101001001110010;
		correct = 32'b00111111101000011001110000110001;
		#400 //-4.384781e-32 * -3.4728764e-32 = 1.2625791
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010110101001111110001000001000;
		b = 32'b01000001000110111110111111111001;
		correct = 32'b00010101000010011100111000101111;
		#400 //2.712295e-25 * 9.746087 = 2.782958e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011110001000001110001010101011;
		b = 32'b00111110000111011010001011001010;
		correct = 32'b10011111100000101010001101111100;
		#400 //-8.517203e-21 * 0.1539413 = -5.5327604e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001100100001000000111110111100;
		b = 32'b11001011011001100110101111101101;
		correct = 32'b01000000100100101011100010100001;
		#400 //-69238240.0 * -15100909.0 = 4.5850377
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110001010000010010011101000011;
		b = 32'b10110010111011100000111100000011;
		correct = 32'b00111101110011111011010111011111;
		#400 //-2.8107514e-09 * -2.7713673e-08 = 0.10142111
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010001000000000011011111111011;
		b = 32'b10110000110111111111001101101000;
		correct = 32'b10011111100100101001000101011100;
		#400 //1.011467e-28 * -1.6294566e-09 = -6.207388e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111111000100001001000110011000;
		b = 32'b11101111000001111100011100011111;
		correct = 32'b11001111100010000100100110001111;
		#400 //1.921648e+38 * -4.20212e+28 = -4573044000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110010110011101001010011100100;
		b = 32'b01011110000000100100000100000000;
		correct = 32'b11010100010010110000000111000110;
		#400 //-8.1835404e+30 * 2.3464458e+18 = -3487632500000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011011000001010001110101100000;
		b = 32'b10111001001000010011100010101110;
		correct = 32'b11100001010100110101111010111011;
		#400 //3.746847e+16 * -0.00015375271 = -2.4369307e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011010011000100111011010101011;
		b = 32'b01111111110101000100100110010110;
		correct = 32'b01111111110101000100100110010110;
		#400 //4.6831564e-23 * nan = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000000001011001101110111011001;
		b = 32'b10100011010100110011101010111110;
		correct = 32'b11011100010100011000000110001100;
		#400 //2.7010405 * -1.1450772e-17 = -2.3588283e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011011011011001001111010111001;
		b = 32'b11001110011011000001001101011001;
		correct = 32'b01001100100000000100101110010010;
		#400 //-6.660261e+16 * -990172740.0 = 67263630.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010101101001010110101111110110;
		b = 32'b11001101001101100001010011101100;
		correct = 32'b10000111111010001001001110100000;
		#400 //6.68133e-26 * -190926530.0 = -3.4994246e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000101100010010011001111011011;
		b = 32'b00010001010110111111011010000101;
		correct = 32'b11110011100111111010111001000111;
		#400 //-4390.482 * 1.7352019e-28 = -2.5302428e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110101001110001111100111101111;
		b = 32'b00010000101100101001011010001001;
		correct = 32'b11100100000001001001010000100101;
		#400 //-6.890904e-07 * 7.0440557e-29 = -9.782581e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111010000100101110100011100000;
		b = 32'b00001110100010110110010111011111;
		correct = 32'b01101011000001101110010111000101;
		#400 //0.0005604159 * 3.4364244e-30 = 1.6308112e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101101000010111000111010101011;
		b = 32'b00111100111101110111000111011100;
		correct = 32'b10101111100100000110000111100101;
		#400 //-7.932914e-12 * 0.03020566 = -2.6263006e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010001011111010010011010101001;
		b = 32'b10001100010111001110100001011111;
		correct = 32'b01000100100100101010111011000011;
		#400 //-1.9970094e-28 * -1.701811e-31 = 1173.4613
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100110001001111111110110001010;
		b = 32'b01110000001010001011000110001110;
		correct = 32'b10110101011111101110111011010001;
		#400 //-1.9832804e+23 * 2.0883253e+29 = -9.49699e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100000001010111100101100101001;
		b = 32'b01110000010110101111110100100110;
		correct = 32'b10101111010010001101010000001011;
		#400 //-4.9516132e+19 * 2.7109508e+29 = -1.8265227e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101011111111011111111010111011;
		b = 32'b00001101001011111101101001101010;
		correct = 32'b01011110001110001110000010111110;
		#400 //1.8047433e-12 * 5.4188945e-31 = 3.3304642e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000011101000001100100011001010;
		b = 32'b00101011000000100111110011101100;
		correct = 32'b01011000000111011011011111111101;
		#400 //321.56866 * 4.635864e-13 = 693654200000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000011000110100101010101110010;
		b = 32'b11010100001000110100100001000000;
		correct = 32'b10101110011100011111100001100100;
		#400 //154.33377 * -2805167300000.0 = -5.501767e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101100010100010001110100001010;
		b = 32'b00000101010110011011101000011000;
		correct = 32'b11100110011101011101111101010101;
		#400 //-2.9716806e-12 * 1.0237471e-35 = -2.9027488e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100010001101111111001100111010;
		b = 32'b11100110011010001100011000000010;
		correct = 32'b10111011010010100100111000010010;
		#400 //8.483201e+20 * -2.748104e+23 = -0.0030869287
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100101110011010110100101100111;
		b = 32'b01011100100011110000010101111001;
		correct = 32'b10001000101101111101011001101010;
		#400 //-3.5633255e-16 * 3.220555e+17 = -1.106432e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101000100001011001001011110111;
		b = 32'b10111100011011000111100111100101;
		correct = 32'b11101011100100001001101000101000;
		#400 //5.046286e+24 * -0.014433359 = -3.496266e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110011010011101111100110110;
		b = 32'b11100100011001111001110111111000;
		correct = 32'b00010001100000010011111100000001;
		#400 //-3.4849631e-06 * -1.7090323e+22 = 2.039144e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001101111000111101101010011111;
		b = 32'b10100110101000111010110110101111;
		correct = 32'b11100110101100100010111111000111;
		#400 //477844450.0 * -1.1357474e-15 = -4.207313e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101111111101100100001100111000;
		b = 32'b00111001101111111110111001011101;
		correct = 32'b01110101101001000011101111100110;
		#400 //1.5242915e+29 * 0.00036607953 = 4.163826e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010111111000110010011110111011;
		b = 32'b00110110111001111101111110010111;
		correct = 32'b10100000011110101100101001110110;
		#400 //-1.4679561e-24 * 6.9103658e-06 = -2.1242812e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011000000010100111010101110010;
		b = 32'b11001010001101100001011101000001;
		correct = 32'b10001101010000101010100001110101;
		#400 //1.7895377e-24 * -2983376.2 = -5.998364e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101100000110110111111011010111;
		b = 32'b10000010011000011100001101111100;
		correct = 32'b01101001001100000101001000100110;
		#400 //-2.2097235e-12 * -1.6586491e-37 = 1.332243e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101100011111111000001100100101;
		b = 32'b00000100010100011110101000000000;
		correct = 32'b11100111100110111100110111111001;
		#400 //-3.631048e-12 * 2.467528e-36 = -1.4715327e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101011101010111001100001001101;
		b = 32'b10111011011100101101110111010101;
		correct = 32'b10101111101101001101111111001111;
		#400 //1.2192553e-12 * -0.0037058492 = -3.2900835e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010100111011010100000111100111;
		b = 32'b11111101100011111010101010100001;
		correct = 32'b00010110110100110110001010010001;
		#400 //-8152103000000.0 * -2.3870695e+37 = 3.4151093e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110100100100111100110100011100;
		b = 32'b01010001000001110101011110110100;
		correct = 32'b01100011000010111100100001100000;
		#400 //9.368015e+31 * 36330750000.0 = 2.578536e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000001010000111110100001011000;
		b = 32'b01111000011011000100010100001100;
		correct = 32'b10001000010101000100010001110000;
		#400 //-12.244225 * 1.9168476e+34 = -6.3876877e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001011001011101110101001100010;
		b = 32'b11011010100100111001101101100000;
		correct = 32'b10110000000101111010111001100001;
		#400 //11463266.0 * -2.077383e+16 = -5.518129e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001001000000000101011010001111;
		b = 32'b01111000101110100011111100010001;
		correct = 32'b10001111101100000110011101011101;
		#400 //-525672.94 * 3.0220199e+34 = -1.7394754e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011001111100100110001101110010;
		b = 32'b10111110001111111101111101010001;
		correct = 32'b00011011001000011011001100101000;
		#400 //-2.5062379e-23 * -0.18737532 = 1.3375496e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110011111110101000110110000000;
		b = 32'b10100110010110011111010111010001;
		correct = 32'b11001101000100110010001111110000;
		#400 //1.1667271e-07 * -7.562014e-16 = -154287870.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001010010100110001100011110111;
		b = 32'b10011101000010011111000100111001;
		correct = 32'b00101100110000111110000111101110;
		#400 //-1.0163976e-32 * -1.8256508e-21 = 5.5673166e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011010110000100010000111110111;
		b = 32'b00101110010000000010110101011101;
		correct = 32'b00101100000000010100110101101101;
		#400 //8.029139e-23 * 4.3696036e-11 = 1.8374983e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001110100010011000110010110011;
		b = 32'b00101011011010111101011111110101;
		correct = 32'b11100010100101010100111000101001;
		#400 //-1153849700.0 * 8.378847e-13 = -1.3770984e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001101101001101110010110101000;
		b = 32'b00110000100110011101100000101111;
		correct = 32'b01011100100010101101110000100011;
		#400 //350008580.0 * 1.1193658e-09 = 3.1268472e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000111011001001011101010101001;
		b = 32'b01101110111010010110110011000000;
		correct = 32'b10010111111110101101100110100111;
		#400 //-58554.66 * 3.612074e+28 = -1.6210815e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100000101111100000001101011000;
		b = 32'b01100101111011011110001110010110;
		correct = 32'b10111010010011000111101010101010;
		#400 //-1.0953507e+20 * 1.4042488e+23 = -0.0007800261
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101010101100010101111100001010;
		b = 32'b01001101100000110101111000101000;
		correct = 32'b11011100101011001101001011110111;
		#400 //-1.0721434e+26 * 275498240.0 = -3.8916523e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111000111011010100101000011111;
		b = 32'b11100111000010110111111010101011;
		correct = 32'b11010001010110011011110001110101;
		#400 //3.8502428e+34 * -6.5874555e+23 = -58448105000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110011101001100100000011100110;
		b = 32'b01000011110111001111100000001011;
		correct = 32'b01101111010000001001110000111111;
		#400 //2.634392e+31 * 441.93784 = 5.961001e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011100110011100110000001100;
		b = 32'b00011100111101110110011101100001;
		correct = 32'b11101110000111110010010000001101;
		#400 //-20158488.0 * 1.6371812e-21 = -1.2312925e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010100001001000111011010010011;
		b = 32'b01010010000111011010101101010100;
		correct = 32'b11000001100001011000001111110111;
		#400 //-2825456000000.0 * 169296070000.0 = -16.689436
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110110111000000001111011011100;
		b = 32'b10111010110010011101011101011111;
		correct = 32'b10111011100011100010000011101111;
		#400 //6.6793127e-06 * -0.0015399269 = -0.004337422
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100100011100110111100011110011;
		b = 32'b01000000111111110000011111001111;
		correct = 32'b11100010111101000110010111100100;
		#400 //-1.7965096e+22 * 7.969703 = -2.2541738e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100111100001110110111100001110;
		b = 32'b01000011011001111000100001100001;
		correct = 32'b11100011100101011011111011101101;
		#400 //-1.2791361e+24 * 231.53273 = -5.524645e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110000011101110010111000101010;
		b = 32'b11101111011110111001111100010110;
		correct = 32'b11000000011110110111101101001011;
		#400 //3.0599443e+29 * -7.787306e+28 = -3.9294002
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100010101100101001101010011100;
		b = 32'b00101111110001110100001011010010;
		correct = 32'b11110010011001010111010111111101;
		#400 //-1.6473306e+21 * 3.6245368e-10 = -4.5449412e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001000001100000100000111001011;
		b = 32'b10001001111101010011100101010111;
		correct = 32'b11111101101110000000000010011011;
		#400 //180487.17 * -5.9035527e-33 = -3.0572637e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010101011111011110000001111011;
		b = 32'b11111100001000111110100111111110;
		correct = 32'b10011000110001100100000001110001;
		#400 //17446286000000.0 * -3.4043613e+36 = -5.124687e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001111011100101111000010000110;
		b = 32'b11001011010110111110100101011100;
		correct = 32'b11000011100011010110011101001011;
		#400 //4075849200.0 * -14412124.0 = -282.80698
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111010011100010011111010100000;
		b = 32'b11001000100100110000111010000111;
		correct = 32'b01110001010100011111101101110111;
		#400 //-3.1315343e+35 * -301172.22 = 1.0397819e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111011101110000100111111000110;
		b = 32'b10011010011010110011111000010010;
		correct = 32'b01100000110010001001001100111000;
		#400 //-0.005624744 * -4.8647e-23 = 1.1562366e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100000111111000100111101011101;
		b = 32'b00010101100110010101100101100001;
		correct = 32'b01001010110100101001101000110001;
		#400 //4.274298e-19 * 6.193722e-26 = 6901016.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101101000001011100101010000101;
		b = 32'b10110100010100010110111011101010;
		correct = 32'b10111000001000111000101000000000;
		#400 //7.605143e-12 * -1.9504992e-07 = -3.899075e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101001100110111010010000011001;
		b = 32'b11100000100011011101111010010100;
		correct = 32'b11001000100011000110110011011100;
		#400 //2.3519804e+25 * -8.178217e+19 = -287590.88
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100001010111001100000100010111;
		b = 32'b10111111011011010101000101000011;
		correct = 32'b10100001011011100010001000000110;
		#400 //7.479445e-19 * -0.9270212 = -8.0682566e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100001110100010011010010110111;
		b = 32'b11011001100110101001010001001100;
		correct = 32'b10000111101011010011101111011011;
		#400 //1.4176344e-18 * -5438775000000000.0 = -2.6065327e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011011100011101110011110100000;
		b = 32'b10101100110101100111011100001011;
		correct = 32'b10101110001010101001010010110011;
		#400 //2.3641614e-22 * -6.0954622e-12 = -3.8785596e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101110111011011101111000100000;
		b = 32'b11001011111010111010001011011111;
		correct = 32'b11100010100000010011011001010000;
		#400 //3.680824e+28 * -30885310.0 = -1.1917718e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100100011101101100011101011000;
		b = 32'b01011101000001110111000111111111;
		correct = 32'b00000110111010010011011010101000;
		#400 //5.3511598e-17 * 6.099914e+17 = 8.772517e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010110001100100111001100001011;
		b = 32'b01000000001101110110001111110001;
		correct = 32'b01010101011110010001101001001011;
		#400 //49051794000000.0 * 2.865475 = 17118208000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001010100110010011100111000011;
		b = 32'b00110000111100111110100100110110;
		correct = 32'b10011001001000001101000111101011;
		#400 //-1.4755092e-32 * 1.774686e-09 = -8.314199e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101010000100110010011111100100;
		b = 32'b10010000001000011100010110010110;
		correct = 32'b11011001011010001101111011011100;
		#400 //1.3070063e-13 * -3.1903866e-29 = -4096702000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011100101100110000110000111;
		b = 32'b01101110111101000000000000101111;
		correct = 32'b10011100000111011100011010111011;
		#400 //-19710734.0 * 3.7757282e+28 = -5.2203796e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111011011110110000010010111101;
		b = 32'b01101001010111000011010001010001;
		correct = 32'b00010001100100011110100101011110;
		#400 //0.0038302385 * 1.6638171e+25 = 2.302079e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010001001100110010101010000100;
		b = 32'b10101101101100101101001100010110;
		correct = 32'b11100011000000000011111010010101;
		#400 //48094527000.0 * -2.0329998e-11 = -2.3656928e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010110110000011101000011101101;
		b = 32'b01011010011000110111011010110001;
		correct = 32'b00111011110110100010000110011001;
		#400 //106551540000000.0 * 1.6006331e+16 = 0.006656837
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110111101100111110001111011000;
		b = 32'b11110100011000001011110000010101;
		correct = 32'b01000010110011001110101010011111;
		#400 //-7.297206e+33 * -7.122127e+31 = 102.458244
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010111010111011001001000010011;
		b = 32'b00100000110101010101011010110001;
		correct = 32'b00110110000001001111000001100110;
		#400 //7.1593323e-25 * 3.614097e-19 = 1.9809463e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110100100101000010000001101001;
		b = 32'b01000011011110111111010010101011;
		correct = 32'b00110000100101101000000100010111;
		#400 //2.759073e-07 * 251.95573 = 1.0950626e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010101110110100010000100100110;
		b = 32'b10100011001100000101001010101111;
		correct = 32'b10110010000111100101100101011010;
		#400 //8.81018e-26 * -9.558488e-18 = -9.217127e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111001000111101101001001000001;
		b = 32'b01000011101100101000101111111100;
		correct = 32'b01110100111000111011011110110101;
		#400 //5.154046e+34 * 357.09363 = 1.4433318e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011010010111100010011101010101;
		b = 32'b01101001111000010001110101101101;
		correct = 32'b10101111111111001010000111100110;
		#400 //-1.5632673e+16 * 3.4018409e+25 = -4.595357e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111001001001111100011100101110;
		b = 32'b11010100110110101101111110001011;
		correct = 32'b01100011110001000011110011011011;
		#400 //-5.444709e+34 * -7520426400000.0 = 7.239894e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101110110011100111101011111110;
		b = 32'b01101101110100010000110001110110;
		correct = 32'b01000000011111001101101011011110;
		#400 //3.19513e+28 * 8.087179e+27 = 3.9508586
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010010111100100001100100001010;
		b = 32'b11101110100011111101011100001001;
		correct = 32'b00100011110101110110111111111101;
		#400 //-519901100000.0 * -2.225816e+28 = 2.3357776e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010111010011010111110000000000;
		b = 32'b00001010110010011001011100011110;
		correct = 32'b01001100000000100111100011111001;
		#400 //6.6395582e-25 * 1.941244e-32 = 34202596.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101100010001000000100000101101;
		b = 32'b01010001100001110110010101101001;
		correct = 32'b11011010001110010101001011010010;
		#400 //-9.479523e+26 * 72690246000.0 = -1.3040983e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001001010000110001101001011111;
		b = 32'b00011111100001110001010100101101;
		correct = 32'b00101001001110001101111110001111;
		#400 //2.348467e-33 * 5.7209756e-20 = 4.1050113e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110010011110010000011110001010;
		b = 32'b11001111000110001110011011110101;
		correct = 32'b01100010110100000111100010111110;
		#400 //-4.9325364e+30 * -2565272800.0 = 1.9228116e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101000010100101100011001010001;
		b = 32'b00101100011000110010111000010111;
		correct = 32'b00111011011011011000001101110010;
		#400 //1.1700345e-14 * 3.2284225e-12 = 0.0036241678
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010110000010011001111010001111;
		b = 32'b10010111101111011101101010101010;
		correct = 32'b11111101101110011001000100000010;
		#400 //37828524000000.0 * -1.2269037e-24 = -3.0832513e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011110010100101100001001001;
		b = 32'b00110010010011011110011111011011;
		correct = 32'b11011000111110111001001010101000;
		#400 //-26521746.0 * 1.1985288e-08 = -2212858400000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010101100111001010111001101000;
		b = 32'b11101010101010100001001011001010;
		correct = 32'b10101010011010111101011101111101;
		#400 //21534110000000.0 * -1.0280306e+26 = -2.0946955e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001000000111101000000111100111;
		b = 32'b01100001100100111101101101001010;
		correct = 32'b10100110000010010011100001110000;
		#400 //-162311.61 * 3.409341e+20 = -4.760791e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110110001110111110111101101101;
		b = 32'b01001111111101000101101100010011;
		correct = 32'b01100101110001001110010000010010;
		#400 //9.52945e+32 * 8199218700.0 = 1.1622387e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011110111001100101010111000101;
		b = 32'b11111011011111100000111010001111;
		correct = 32'b00100010111010000001100011000100;
		#400 //-8.2986943e+18 * -1.3191387e+36 = 6.2909948e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111111101111011110100100001111;
		b = 32'b10111010001000010100011000110010;
		correct = 32'b01000101000101101011101001011011;
		#400 //-1.4836749 * -0.00061521225 = 2411.6472
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001011000011001101110011101100;
		b = 32'b00110010010000001010011001001001;
		correct = 32'b01011000001110110010111100011101;
		#400 //9231596.0 * 1.121368e-08 = 823244100000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010011101000110010000110001010;
		b = 32'b11000000010001100110100000000001;
		correct = 32'b00010010110100100111110000101000;
		#400 //-4.1180057e-27 * -3.100098 = 1.328347e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010100111111100000011100101110;
		b = 32'b10100010001000011111110010101100;
		correct = 32'b10110010010010001011101011001001;
		#400 //2.5650278e-26 * -2.1953332e-18 = -1.1684002e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100011010101001110101101000101;
		b = 32'b11110010101110111111011011111010;
		correct = 32'b00110000000100001111111001001011;
		#400 //-3.9276627e+21 * -7.446051e+30 = 5.2748267e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001100000110001010101000000100;
		b = 32'b01011001110101111101101001101011;
		correct = 32'b00110001101101010000111011101110;
		#400 //40019984.0 * 7594659000000000.0 = 5.2694906e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100100100101011111001010100001;
		b = 32'b00010111100111111010010110110111;
		correct = 32'b01001100011100000111001001001001;
		#400 //6.502948e-17 * 1.0316966e-24 = 63031588.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011100000101100001000000001010;
		b = 32'b00010011001101110101111100010010;
		correct = 32'b01001000010100010111111110100010;
		#400 //4.9651567e-22 * 2.314472e-27 = 214526.53
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111110101100110100010110110011;
		b = 32'b00000101111001101100100001011101;
		correct = 32'b11111000010001101101110001110010;
		#400 //-0.35014114 * 2.1702698e-35 = -1.613353e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010100110111111010111001011001;
		b = 32'b01001100011011001010001101001110;
		correct = 32'b01000111111100011111101110100101;
		#400 //7685622000000.0 * 62033210.0 = 123895.29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100100100100000011100010000011;
		b = 32'b00110000011010100010111111011111;
		correct = 32'b10110011100111011010011101101011;
		#400 //-6.254578e-17 * 8.5196733e-10 = -7.3413354e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000000110100101101000001110010;
		b = 32'b11100000100100101101001000111000;
		correct = 32'b00011111101101111100101000101100;
		#400 //-6.587945 * -8.463664e+19 = 7.783798e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001001011001010101010000101010;
		b = 32'b00111110110011010000010011101110;
		correct = 32'b10001010000011110010110101011101;
		#400 //-2.7604446e-33 * 0.40042824 = -6.8937314e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100000111000101001011101011110;
		b = 32'b10110110010101110101001000110100;
		correct = 32'b00101010000001101011001100011110;
		#400 //-3.8386056e-19 * -3.2085345e-06 = 1.1963735e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011111001101110010101100001111;
		b = 32'b00101101010010101100110010111011;
		correct = 32'b00110001011001110011011111110011;
		#400 //3.8787375e-20 * 1.152783e-11 = 3.3646728e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001100110001101101001100001001;
		b = 32'b11110011010110110100110011100100;
		correct = 32'b10011000111010000001100011101101;
		#400 //104241224.0 * -1.7374764e+31 = -5.9995763e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000000000111001110110000111111;
		b = 32'b11001100110010101010111101111111;
		correct = 32'b00110010110001100011001100101011;
		#400 //-2.4519193 * -106265590.0 = 2.3073502e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000011010010111111101100111010;
		b = 32'b11100100110111110101000001001110;
		correct = 32'b00011101111010011101011010000111;
		#400 //-203.98135 * -3.2955284e+22 = 6.1896403e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001101101111001010011101000011;
		b = 32'b00101001100101000011111001011001;
		correct = 32'b11100011101000101110010001000001;
		#400 //-395634780.0 * 6.583336e-14 = -6.00964e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001011010110100011111100000111;
		b = 32'b11111111111101100100001000100110;
		correct = 32'b11111111111101100100001000100110;
		#400 //-4.203269e-32 * nan = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001010011000110011011001111111;
		b = 32'b01111101101011010100011000000111;
		correct = 32'b00001100001001111101100010001011;
		#400 //3722655.8 * 2.8790006e+37 = 1.2930376e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000011001111001001110001000111;
		b = 32'b10001110010101100110001010010110;
		correct = 32'b10110100011000010011100011100000;
		#400 //5.542763e-37 * -2.6425004e-30 = -2.0975449e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010100110011110011011001110111;
		b = 32'b10110000110010001100010000110111;
		correct = 32'b01100011100001000001110000100001;
		#400 //-7119776000000.0 * -1.4607683e-09 = 4.873994e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111100100100000110101101000111;
		b = 32'b11010101110000011101011111010101;
		correct = 32'b00100110001111101011101001010101;
		#400 //-0.017629279 * -26641592000000.0 = 6.617202e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010011110011110100110110010011;
		b = 32'b11101010011110100010100110110110;
		correct = 32'b00101000110101000010001111011010;
		#400 //-1780719400000.0 * -7.5607107e+25 = 2.3552276e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101001011001100001000110011110;
		b = 32'b00101100100110001010000001010011;
		correct = 32'b11111100010000001111001001111011;
		#400 //-1.7383508e+25 * 4.3378994e-12 = -4.0073563e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000110101111100001000011110101;
		b = 32'b10011000010110110101110110111100;
		correct = 32'b10101101110111011100111010011010;
		#400 //7.149497e-35 * -2.835241e-24 = -2.521654e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111010011100000111000011111111;
		b = 32'b11100100111111100110110011110111;
		correct = 32'b01010100111100011110110111100001;
		#400 //-3.1211077e+35 * -3.7546598e+22 = 8312624500000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001100100101101100101000011101;
		b = 32'b00000011100000100000101110101100;
		correct = 32'b11001000100101000110101011101001;
		#400 //-2.3232802e-31 * 7.643393e-37 = -303959.28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101110101100110110101001100110;
		b = 32'b01010001111100001000111100011101;
		correct = 32'b01011100001111101110111010010010;
		#400 //2.7763222e+28 * 129149150000.0 = 2.1497023e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111010101011101101011011101101;
		b = 32'b11101101001010110110110000000010;
		correct = 32'b10001101000000101000110101001100;
		#400 //0.0013339199 * -3.315782e+27 = -4.0229423e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001111001011110111101010101010;
		b = 32'b00100000101010001101001001110010;
		correct = 32'b01101110000001010000110000100001;
		#400 //2944051700.0 * 2.8599568e-19 = 1.0294042e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101000100110110001010000110100;
		b = 32'b11000001100110111100011110110010;
		correct = 32'b11100110011111101101100100001000;
		#400 //5.858716e+24 * -19.472507 = -3.0087115e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110000100101110111111011000001;
		b = 32'b11101100111001110110011000011110;
		correct = 32'b10000011001001111001100111101110;
		#400 //1.1022722e-09 * -2.2379528e+27 = -4.925359e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111100000101111011001001101110;
		b = 32'b01010100110000110000001000001010;
		correct = 32'b10100110110001110010010010001110;
		#400 //-0.00925885 * 6700422700000.0 = -1.3818307e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111001110000110000011010011111;
		b = 32'b00111001011011111001100010111111;
		correct = 32'b10111111110100000110000010110110;
		#400 //-0.0003719823 * 0.00022849719 = -1.6279514
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100011011010010100010101000110;
		b = 32'b10100100110001001001110101101101;
		correct = 32'b10111110000101111101110100001111;
		#400 //1.26456245e-17 * -8.526814e-17 = -0.14830421
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010101001111100000010101000110;
		b = 32'b01010011011010000101100110011010;
		correct = 32'b01000001010100010101110010101111;
		#400 //13058116000000.0 * 997935700000.0 = 13.085128
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110011000001111111111101001000;
		b = 32'b10001011101011100001100100101111;
		correct = 32'b11100110110001111111100110001010;
		#400 //3.1664314e-08 * -6.7060254e-32 = -4.7217706e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111100100001100101011011000001;
		b = 32'b00100101010110111110111100111011;
		correct = 32'b11010110100111000101111001000000;
		#400 //-0.01639879 * 1.9076276e-16 = -85964310000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000001101011111100010001101101;
		b = 32'b10010010000000010110110100001111;
		correct = 32'b01101111001011011101010010101000;
		#400 //-21.970911 * -4.083965e-28 = 5.379799e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000010110111000000110111100111;
		b = 32'b11010010101100010011111011011000;
		correct = 32'b00101111100111101110101000111000;
		#400 //-110.02715 * -380631780000.0 = 2.8906455e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011101111000011010010010011001;
		b = 32'b10100001110100001010011100011101;
		correct = 32'b00111011100010100110110000111011;
		#400 //-5.9727194e-21 * -1.4138863e-18 = 0.004224328
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110110010010011111100001101;
		b = 32'b10111001000011101000011101011101;
		correct = 32'b00111101001101001011101101101100;
		#400 //-5.997607e-06 * -0.00013592602 = 0.044124052
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001111010010110100110001100111;
		b = 32'b10001011100000011011010011010001;
		correct = 32'b11000011010010001001111110111111;
		#400 //1.0023387e-29 * -4.9961055e-32 = -200.62401
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001000110000100000110011110011;
		b = 32'b11101110010110011110101000111011;
		correct = 32'b10011001111000111111011100000000;
		#400 //397415.6 * -1.6860354e+28 = -2.3571012e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110001110110001110011101000010;
		b = 32'b00010001101001011001000111001000;
		correct = 32'b01011111101001111010111110001001;
		#400 //6.3127183e-09 * 2.6122255e-28 = 2.4166054e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011000111101110001100001001111;
		b = 32'b00011111011011100011001000111000;
		correct = 32'b00111001000001001100100000101111;
		#400 //6.387255e-24 * 5.044e-20 = 0.00012663075
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010110001110000111110011100110;
		b = 32'b01000011110001000010110011001110;
		correct = 32'b00010001111100001011111110110001;
		#400 //1.4902813e-25 * 392.35004 = 3.7983462e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101001000011000011110010000000;
		b = 32'b10000100101111000100010111111111;
		correct = 32'b11100011101111101010111011001011;
		#400 //3.113872e-14 * -4.426287e-36 = -7.034953e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111011000001001011000101110001;
		b = 32'b11101101110110110001010101100101;
		correct = 32'b11001100100110110000110101101100;
		#400 //6.889821e+35 * -8.475385e+27 = -81292130.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000001101110011000111010000001;
		b = 32'b10011110010000001011100100111110;
		correct = 32'b00100010111101100111101011011110;
		#400 //-6.816275e-38 * -1.02027026e-20 = 6.6808524e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001110100000110110100100011000;
		b = 32'b11100110110100110001111100011101;
		correct = 32'b10100111000111110101100000111101;
		#400 //1102351400.0 * -4.9849663e+23 = -2.2113517e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101111000101001111010010001011;
		b = 32'b01010111101100101001011000100111;
		correct = 32'b11010110110101011000011000110001;
		#400 //-4.6099416e+28 * 392715940000000.0 = -117386160000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111010100000100111000010011;
		b = 32'b01100101111010001010010101111100;
		correct = 32'b10010000111001010011011100010001;
		#400 //-1.2415944e-05 * 1.3733021e+23 = -9.0409417e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100111010101000010010110011111;
		b = 32'b10101110101101101000001100011001;
		correct = 32'b10111000000101001100100010011011;
		#400 //2.9441305e-15 * -8.2996894e-11 = -3.5472778e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000100100000111110110001010010;
		b = 32'b00101001011011001100110110000111;
		correct = 32'b10011010100011101001111000101110;
		#400 //-3.1014978e-36 * 5.2580793e-14 = -5.8985377e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011011011100001101010011111;
		b = 32'b11101011100101100010111110000010;
		correct = 32'b00011111010010101110111001010111;
		#400 //-15604383.0 * -3.6312644e+26 = 4.2972314e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001100001000100101100011001101;
		b = 32'b10000111111111001111100101101000;
		correct = 32'b11000011101001000100100111100110;
		#400 //1.2506749e-31 * -3.8063334e-34 = -328.57733
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001001110011101110101011110001;
		b = 32'b01001011011100101001101100101100;
		correct = 32'b00111101110110100101011101100000;
		#400 //1695070.1 * 15899436.0 = 0.10661197
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010111011101000110010001001101;
		b = 32'b01001000000001100000000000010100;
		correct = 32'b00001110111010010111001011000111;
		#400 //7.896725e-25 * 137216.31 = 5.754946e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010000110111100111100001010010;
		b = 32'b10100000001000011010010101110010;
		correct = 32'b01110000001100000010100111010110;
		#400 //-29859418000.0 * -1.3691972e-19 = 2.1807975e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110110110110110111101010001010;
		b = 32'b11111001110101010100010010001001;
		correct = 32'b10111100100000111011101001001100;
		#400 //2.2257781e+33 * -1.3841866e+35 = -0.016080044
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011000001001110110100000011101;
		b = 32'b10101000101101011101111011001101;
		correct = 32'b01101110111010111010010000011100;
		#400 //-736262400000000.0 * -2.0191661e-14 = 3.6463687e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011010100011010001111101101010;
		b = 32'b11001011011101010000111101110000;
		correct = 32'b01001110100100110110110000101100;
		#400 //-1.9861256e+16 * -16060272.0 = 1236670000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010010110011011110011101011000;
		b = 32'b10010110110011110101110100110011;
		correct = 32'b11111011011111100011001001110110;
		#400 //442174800000.0 * -3.350147e-25 = -1.3198669e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111111001110001011011100101000;
		b = 32'b11101000101011010111001111000010;
		correct = 32'b00010110000010000100111111010010;
		#400 //-0.72154474 * -6.552838e+24 = 1.1011179e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100010111111101101010100100111;
		b = 32'b00101100011000010100101001111010;
		correct = 32'b11110110000100001100100011000100;
		#400 //-2.3504161e+21 * 3.2015766e-12 = -7.341433e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010100000101101101000110101101;
		b = 32'b10111110010001000000100001000011;
		correct = 32'b00010101010001001111010010101010;
		#400 //-7.614416e-27 * -0.19143777 = 3.977489e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110111110011110110110101000011;
		b = 32'b01100110000101100101001101110011;
		correct = 32'b01010001001100001001111011010001;
		#400 //8.414231e+33 * 1.7747358e+23 = 47411170000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000011100101011011000010101;
		b = 32'b10010101110111011100001010110100;
		correct = 32'b01011010000011000001011110111101;
		#400 //-8.829784e-10 * -8.9568377e-26 = 9858149000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011111010011111001111011011000;
		b = 32'b00100001110100100110011011000001;
		correct = 32'b00111100111111001001110111001110;
		#400 //4.3965347e-20 * 1.4257352e-18 = 0.030836966
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011101100111111010111001011011;
		b = 32'b00011101110110001000111011011100;
		correct = 32'b10111111001111001100001110010011;
		#400 //-4.226723e-21 * 5.7322437e-21 = -0.7373592
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010010111101000001111101100000;
		b = 32'b00001001100010111001010011001001;
		correct = 32'b11001000110111111101111000010010;
		#400 //-1.5406299e-27 * 3.360295e-33 = -458480.56
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001111010001110101110001110000;
		b = 32'b10001010111011010111011000100111;
		correct = 32'b01000011110101101110110011010010;
		#400 //-9.82926e-30 * -2.2866714e-32 = 429.85016
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110010011110111101110010101100;
		b = 32'b10111101101000000110110100111011;
		correct = 32'b00110100010010001111010000100110;
		#400 //-1.4660298e-08 * -0.07833334 = 1.8715272e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000111111010010001100111001;
		b = 32'b10100011100100111100110011010101;
		correct = 32'b01001100110110110011100111010011;
		#400 //-1.8418184e-09 * -1.6024522e-17 = 114937496.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100111010011100110010011001000;
		b = 32'b01110001010111111111110111110101;
		correct = 32'b10110101011010111110001100001011;
		#400 //-9.746666e+23 * 1.10915476e+30 = -8.7874713e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011100100011100000000010000011;
		b = 32'b01000111110011111011010110111110;
		correct = 32'b00010100001011110000010000001001;
		#400 //9.396904e-22 * 106347.484 = 8.836038e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110000000110100011000100000010;
		b = 32'b00010011110100110000001110010100;
		correct = 32'b01011011101110110001000001000000;
		#400 //5.609452e-10 * 5.3267417e-27 = 1.05307375e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111111011101111101110110110001;
		b = 32'b01110000011010101101011110101010;
		correct = 32'b00001110100001110001100100110011;
		#400 //0.9682265 * 2.9072086e+29 = 3.3304335e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101000101110001100100111011111;
		b = 32'b10011101011000011000100110011101;
		correct = 32'b01001010110100011011111101001001;
		#400 //-2.0515651e-14 * -2.9849646e-21 = 6872996.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001100101110110001110001010110;
		b = 32'b11100000110110101010000000110111;
		correct = 32'b00101011010110110001100011101010;
		#400 //-98099890.0 * -1.2602922e+20 = 7.7839005e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101000110001111001001110111100;
		b = 32'b00101011110011111000110101100110;
		correct = 32'b10111100011101100010100111000011;
		#400 //-2.2157508e-14 * 1.4747481e-12 = -0.015024605
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111011001010110111101011011001;
		b = 32'b00010110101000100011100101101111;
		correct = 32'b11100100000001110100110110001010;
		#400 //-0.0026165752 * 2.6208757e-25 = -9.983591e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011101110110100101101111100;
		b = 32'b11010000100000111010111101110100;
		correct = 32'b00111010101101100000110110011111;
		#400 //-24549112.0 * -17674510000.0 = 0.0013889557
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000110000001001010001010010000;
		b = 32'b10010110100111101010111001001000;
		correct = 32'b10101110110101011111101011110101;
		#400 //2.4945873e-35 * -2.5636264e-25 = -9.7306975e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100011010011011110100100110100;
		b = 32'b01000100110110101110011011110001;
		correct = 32'b10011101111100001100111010100100;
		#400 //-1.1162455e-17 * 1751.2169 = -6.3741132e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100101100000110010101100011010;
		b = 32'b10001101010111101100100000111010;
		correct = 32'b11010111100101101011100111100111;
		#400 //2.2754084e-16 * -6.8650046e-31 = -331450380000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101110110011111111001110000100;
		b = 32'b00111100011001111101000010100101;
		correct = 32'b01110001111001011010010110000011;
		#400 //3.2178895e+28 * 0.014148866 = 2.2743091e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100011100111011000111110110111;
		b = 32'b11010000111101000011010011010101;
		correct = 32'b00010010001001010010101110101101;
		#400 //-1.708284e-17 * -32776825000.0 = 5.2118654e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001111101100010011011011001110;
		b = 32'b01000100100000000111010110010001;
		correct = 32'b10001010101100001001010010011110;
		#400 //-1.7474658e-29 * 1027.674 = -1.7004087e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100111000101101100001001100001;
		b = 32'b11001101010001100001010010110000;
		correct = 32'b11011001010000101101011101110010;
		#400 //7.119406e+23 * -207702780.0 = -3427689400000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000010000100001111111010000;
		b = 32'b01001000111100100111011001001001;
		correct = 32'b10100110110011001111011010011000;
		#400 //-7.0621997e-10 * 496562.28 = -1.4222183e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100100110011010111000010001101;
		b = 32'b10111010010111010111110011011110;
		correct = 32'b01101001111011010111001110000111;
		#400 //-3.0317541e+22 * -0.00084490876 = 3.5882623e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100000010100110100010100001111;
		b = 32'b00101010100011001101010001100100;
		correct = 32'b00110101010000000000010111100010;
		#400 //1.7895245e-19 * 2.501637e-13 = 7.1534134e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011000110111010110011110101011;
		b = 32'b01010000100010001100010100100000;
		correct = 32'b01000111110011110011010100111100;
		#400 //1947498600000000.0 * 18356961000.0 = 106090.47
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011001011101001000111010011010;
		b = 32'b01000010010000000101101101001010;
		correct = 32'b00010110101000101011110001011100;
		#400 //1.26433025e-23 * 48.08915 = 2.6291383e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000010001010100010100010101011;
		b = 32'b10001010001101101100000010010111;
		correct = 32'b01110111011011100101101111101100;
		#400 //-42.539715 * -8.7992034e-33 = 4.8344963e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001001110010110111000101000111;
		b = 32'b00111010101010000001100010010010;
		correct = 32'b10001110100110101110101001010001;
		#400 //-4.8976998e-33 * 0.0012824705 = -3.818957e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100111110000100000011100010011;
		b = 32'b01011110001011001111011000110100;
		correct = 32'b01001001000011111001011011111100;
		#400 //1.8325392e+24 * 3.1158015e+18 = 588143.75
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011101110100100000001010110111;
		b = 32'b11000000111000110011010100111011;
		correct = 32'b00011100011011001001111110011000;
		#400 //-5.5589344e-21 * -7.100248 = 7.829212e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111111001000101000001101101111;
		b = 32'b01111110100101101011001010001100;
		correct = 32'b11000000000010100000100101001010;
		#400 //-2.1601738e+38 * 1.0015563e+38 = -2.156817
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000110011110001011000010000110;
		b = 32'b00101010100000011001001100111110;
		correct = 32'b10011011011101011010101010011000;
		#400 //-4.6773305e-35 * 2.3017173e-13 = -2.0321047e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000110100000010010110011100100;
		b = 32'b00001001011101101000010100100000;
		correct = 32'b10111100100001100010010010010000;
		#400 //-4.859037e-35 * 2.9673768e-33 = -0.016374856
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000110111010101101001111000010;
		b = 32'b10001000010111100110101111001110;
		correct = 32'b10111110000001110010001110110111;
		#400 //8.8332167e-35 * -6.693242e-34 = -0.13197218
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111000101010001010000001011001;
		b = 32'b00001110100100011101000101111110;
		correct = 32'b01101001100101000000010101100000;
		#400 //8.040731e-05 * 3.5946993e-30 = 2.23683e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111001000010111101110101100;
		b = 32'b11011100110110000010101010000101;
		correct = 32'b10101001101111110011110110000101;
		#400 //41339.67 * -4.8676277e+17 = -8.492776e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000100110110010011000001100011;
		b = 32'b00011110001000110000000001010011;
		correct = 32'b10100110001010101000110101010000;
		#400 //-5.106089e-36 * 8.629215e-21 = -5.917211e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011101000110111010101111000000;
		b = 32'b00001100001100111111010000000111;
		correct = 32'b11010000010111010111010011000110;
		#400 //-2.0602872e-21 * 1.3863093e-31 = -14861670000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011111111000101110011111101011;
		b = 32'b10011101101111100011111000001100;
		correct = 32'b01000001100110001010101100001111;
		#400 //-9.60984e-20 * -5.0356736e-21 = 19.083525
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001101111111111011111100101001;
		b = 32'b00101101111111101001000100111110;
		correct = 32'b10011111100000001001011111001111;
		#400 //-1.57616085e-30 * 2.8940957e-11 = -5.4461255e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110100010110010001011001010111;
		b = 32'b01011110011010110011011110001001;
		correct = 32'b10010101011011000100010010111001;
		#400 //-2.0217827e-07 * 4.2372916e+18 = -4.7714033e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111010010111101101110101111101;
		b = 32'b11100010001111100111000011001101;
		correct = 32'b11010111100101011100101100011011;
		#400 //2.8929555e+35 * -8.782524e+20 = -329399130000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110111101100100111100001101010;
		b = 32'b11001011010000111001001111100100;
		correct = 32'b10101011111010011001101110000100;
		#400 //2.1275326e-05 * -12817380.0 = -1.659881e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011010011011001101111001001011;
		b = 32'b00100001100000101111101011011110;
		correct = 32'b10111000011001110111101010110011;
		#400 //-4.8983223e-23 * 8.875547e-19 = -5.5188964e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010110101100010000000101100100;
		b = 32'b01111000011010001110010100100000;
		correct = 32'b00011101110000101001000011010100;
		#400 //97309765000000.0 * 1.8894689e+34 = 5.150112e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101101001010000101011000000001;
		b = 32'b11001100111000110111110100111111;
		correct = 32'b01011111101111010110111011100011;
		#400 //-3.256091e+27 * -119269880.0 = 2.7300194e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100111100001000010111001011001;
		b = 32'b11000001001110111110110100000110;
		correct = 32'b10100101101101000000111111101101;
		#400 //3.668761e-15 * -11.745367 = -3.1235814e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000111000111101001001110111110;
		b = 32'b11000100101111100111100110010001;
		correct = 32'b01000001110101010010000100001110;
		#400 //-40595.742 * -1523.799 = 26.64114
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110000010000010010101010101111;
		b = 32'b00110111111101111110111111000100;
		correct = 32'b01110111110001110111001011101100;
		#400 //2.3912883e+29 * 2.9556344e-05 = 8.090609e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111001010111010011101101101001;
		b = 32'b01010000111101011111001101101100;
		correct = 32'b01100111111001100100010101110000;
		#400 //7.179391e+34 * 33010967000.0 = 2.1748504e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001000100001000111111111101010;
		b = 32'b10001111010011000101111011101101;
		correct = 32'b10111000101001011111100011110000;
		#400 //7.9745335e-34 * -1.00762586e-29 = -7.914181e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100100011101111111111111011001;
		b = 32'b11111110011100100001000110111100;
		correct = 32'b10100101100000110010001010111101;
		#400 //1.8299126e+22 * -8.0441314e+37 = -2.2748417e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011110111110000100001101100011;
		b = 32'b10101010111001011100110011011111;
		correct = 32'b01110011100010100100100010110010;
		#400 //-8.9446255e+18 * -4.082073e-13 = 2.191197e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110011101100101110000001011001;
		b = 32'b11010011110111111010000101001001;
		correct = 32'b11011111010011001100010010110010;
		#400 //2.834409e+31 * -1920967200000.0 = -1.4755114e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100100111101000111111100111001;
		b = 32'b11011101100011000100101000100010;
		correct = 32'b01000110110111110001010000100011;
		#400 //-3.6081383e+22 * -1.2636162e+18 = 28554.068
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000110101000111100010001110110;
		b = 32'b10110111100011110010011000100100;
		correct = 32'b10001110100100100110111110111100;
		#400 //6.160246e-35 * -1.7064689e-05 = -3.6099375e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100001101110100010101001000110;
		b = 32'b01000111011010100100110111000111;
		correct = 32'b11011001110010110110011101011100;
		#400 //-4.2926756e+20 * 59981.777 = -7156633000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110100101110101010001100001100;
		b = 32'b01011000101010011010000000001100;
		correct = 32'b11011011100011001101011001001110;
		#400 //-1.1829519e+32 * 1492038900000000.0 = -7.9284254e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100110110101011000000110100011;
		b = 32'b01010110011010000101010111110000;
		correct = 32'b00001111111010110100000010111100;
		#400 //1.4814982e-15 * 63863950000000.0 = 2.3197724e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000011010011101101011100000010;
		b = 32'b01111011110011010100001001110000;
		correct = 32'b00000111000000001111110001001010;
		#400 //206.83987 * 2.1315367e+36 = 9.703791e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000001010110101111110011101000;
		b = 32'b00101010001110010011101001010011;
		correct = 32'b10010110100101110101010001100001;
		#400 //-4.0221728e-38 * 1.6451536e-13 = -2.4448616e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110010100010000110011101101100;
		b = 32'b10110101100101100100111001101011;
		correct = 32'b00111100011010000101001001011100;
		#400 //-1.5879515e-08 * -1.1198694e-06 = 0.014179792
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011000110110001110111101011111;
		b = 32'b11100111100111001000111111111010;
		correct = 32'b00110000101100010101101111001100;
		#400 //-1908180800000000.0 * -1.4786901e+24 = 1.2904535e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101010101000000001111011011101;
		b = 32'b10100001000110010011001010111110;
		correct = 32'b01001001000001011100100010100100;
		#400 //-2.8443125e-13 * -5.1905573e-19 = 547978.25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111001111111011110100110101001;
		b = 32'b10110111011011110100111001011100;
		correct = 32'b01000010000001111101000000010100;
		#400 //-0.0004843001 * -1.4263755e-05 = 33.9532
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011001001000100110101000000;
		b = 32'b01000010000000010110100110101000;
		correct = 32'b11001000101000101000001000011000;
		#400 //-10767680.0 * 32.35318 = -332816.75
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010010110101110011111101000110;
		b = 32'b00111101000010001010001000100101;
		correct = 32'b00010101010010011010010101111110;
		#400 //1.3584006e-27 * 0.033357758 = 4.0722177e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110110011010101111010001010011;
		b = 32'b01100011110000010101110000000001;
		correct = 32'b11010010000110111000100011111001;
		#400 //-1.1913603e+33 * 7.1337024e+21 = -167004490000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011011101010011011011001100000;
		b = 32'b01001100100010011110010001111110;
		correct = 32'b01001110100111011000100101111101;
		#400 //9.553959e+16 * 72295410.0 = 1321516700.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010011101010111010011001101011;
		b = 32'b11010000011100001101011000000100;
		correct = 32'b11000010101101100111010100110110;
		#400 //1474462900000.0 * -16162230000.0 = -91.22893
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110101100011100110000110011111;
		b = 32'b11011100101011111111101110101001;
		correct = 32'b11011000010011110001111010111101;
		#400 //3.6097956e+32 * -3.962786e+17 = -910923700000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111000101100011110101000000000;
		b = 32'b01100100100100000010110110101001;
		correct = 32'b01010011100111011111001101000000;
		#400 //2.8868207e+34 * 2.127697e+22 = 1356781800000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000001000100010100110101110111;
		b = 32'b11011011111001101111110111111011;
		correct = 32'b10100100101000010000100010010011;
		#400 //9.081412 * -1.30037e+17 = -6.9837145e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010110011011010110001100001110;
		b = 32'b10010011010111100011100000011011;
		correct = 32'b01000010100010001011110010011100;
		#400 //-1.9175964e-25 * -2.8048001e-27 = 68.36838
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110011101101000101011111010100;
		b = 32'b00010011111011000111101100011110;
		correct = 32'b01011111010000110011101010000010;
		#400 //8.397879e-08 * 5.969618e-27 = 1.4067699e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110011100000010001111010101100;
		b = 32'b11011111110100100111110100111001;
		correct = 32'b01010011000111010000100110010100;
		#400 //-2.045985e+31 * -3.0334684e+19 = 674470560000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011110000101111101000010010100;
		b = 32'b01010010110111010010111100010111;
		correct = 32'b11001010101011111011011000101001;
		#400 //-2.7348516e+18 * 474988900000.0 = -5757716.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101011001000000110011101101000;
		b = 32'b01000100000010101110111000100010;
		correct = 32'b10100110100100111100100011001000;
		#400 //-5.6986924e-13 * 555.7208 = -1.0254596e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001000100001110111101110100011;
		b = 32'b00001000100110101001010010011110;
		correct = 32'b00111111011000000101111101100011;
		#400 //8.154084e-34 * 9.303478e-34 = 0.8764555
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100110100101000100111001100101;
		b = 32'b00111100011111110001010110011101;
		correct = 32'b10101001100101001101011010101011;
		#400 //-1.0290812e-15 * 0.015569118 = -6.609759e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000001010101010100000100110101;
		b = 32'b00011010010101000011001101010010;
		correct = 32'b10100110100000001010001011001100;
		#400 //-3.9168705e-38 * 4.388203e-23 = -8.92591e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001010100001001011001111001000;
		b = 32'b11111011001001010000010101110000;
		correct = 32'b10001110110011011101110011110011;
		#400 //4348388.0 * -8.568393e+35 = -5.0749168e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100110111000111000010011110101;
		b = 32'b11011000001010111111100001010011;
		correct = 32'b01001110001010010101100010100100;
		#400 //-5.372149e+23 * -756332100000000.0 = 710289660.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001101100101011100010111100110;
		b = 32'b10111010110010001001000001101100;
		correct = 32'b10010010001111110010101110010110;
		#400 //9.230476e-31 * -0.001530183 = -6.0322697e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101111100000111110110111000111;
		b = 32'b01010111100101011110011010001111;
		correct = 32'b11010111011000010100111011001011;
		#400 //-8.165998e+28 * 329634950000000.0 = -247728530000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010111010000111111111110011111;
		b = 32'b11000101011010000100100111100000;
		correct = 32'b00010001010110000000000101101100;
		#400 //-6.3330537e-25 * -3716.6172 = 1.7039834e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011001000110011110100000001100;
		b = 32'b01000101010000110001001111101110;
		correct = 32'b11010011010010011111100010001100;
		#400 //-2707550600000000.0 * 3121.2456 = -867458350000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001000000001000100001100001010;
		b = 32'b00010011010010010101010010000100;
		correct = 32'b10110100001010000010110100111100;
		#400 //-3.980111e-34 * 2.5411436e-27 = -1.5662675e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010000111000010111001000100101;
		b = 32'b00000010101001010001001010110011;
		correct = 32'b11001101101011101101000001100000;
		#400 //-8.892272e-29 * 2.4255304e-37 = -366611460.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011011001110101001111011110100;
		b = 32'b11001100100011101100110000001101;
		correct = 32'b00001110001001110100100001011101;
		#400 //-1.543692e-22 * -74866790.0 = 2.061918e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101111111111101001110010000111;
		b = 32'b10110101111011010010100111000101;
		correct = 32'b11111001100010010110101011000100;
		#400 //1.57596845e+29 * -1.7670033e-06 = -8.918877e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110000010000000111100001111101;
		b = 32'b11111010011101001001110101011000;
		correct = 32'b00110101010010010110110111010101;
		#400 //-2.3826713e+29 * -3.1752794e+35 = 7.503816e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101000111011101100000001010001;
		b = 32'b00001101001110111000100000010110;
		correct = 32'b11011011001000101111010111000110;
		#400 //-2.6506712e-14 * 5.778763e-31 = -4.5869177e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011111010101001101111001010110;
		b = 32'b10111010010111001010101100110101;
		correct = 32'b10100100011101101111001101101001;
		#400 //4.5076658e-20 * -0.0008417846 = -5.3548923e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001110011111010001011100010000;
		b = 32'b10111110100111011110100100001110;
		correct = 32'b10001111010011010010011011000001;
		#400 //3.1195762e-30 * -0.3084187 = -1.0114744e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110111111010110110001011001111;
		b = 32'b11101101001110011000110100111101;
		correct = 32'b11001010001000100110000010011101;
		#400 //9.5483894e+33 * -3.589092e+27 = -2660391.2
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101000111011101011110110110111;
		b = 32'b10101100010100101101000111110011;
		correct = 32'b10111100000100001111001111001001;
		#400 //2.6505584e-14 * -2.995934e-12 = -0.008847185
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100100010010010101001011110101;
		b = 32'b00110101010110101101100110111000;
		correct = 32'b00101110011010110111111110011110;
		#400 //4.3655195e-17 * 8.152815e-07 = 5.354616e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001110011111101101010111100111;
		b = 32'b11100110010010101100011111001111;
		correct = 32'b10100111101000001101101111000001;
		#400 //1068857800.0 * -2.3940096e+23 = -4.464718e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001110100010110111000110011100;
		b = 32'b01011011001010111010001010110101;
		correct = 32'b00110010110011111111110000100011;
		#400 //1169739300.0 * 4.831112e+16 = 2.421263e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011000010100101100010101000111;
		b = 32'b01000110111001111110100110111010;
		correct = 32'b00010000111010001010100101100111;
		#400 //2.7241463e-24 * 29684.863 = 9.176887e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100100010110011001011011100001;
		b = 32'b11100011111111011011110101110001;
		correct = 32'b10111111110110111000011100000010;
		#400 //1.6055262e+22 * -9.361354e+21 = -1.7150576
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101011101101110110011000111110;
		b = 32'b01000100101110100111001001010010;
		correct = 32'b01100110011110111101000011101010;
		#400 //4.434325e+26 * 1491.5725 = 2.9729194e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011101110000101001111111100001;
		b = 32'b00001110101000010011101010101110;
		correct = 32'b11001110100110101000001100110111;
		#400 //-5.1516683e-21 * 3.974607e-30 = -1296145300.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010010000011001010000001111000;
		b = 32'b01100001011011010000101110100100;
		correct = 32'b00110000000101111101111100011111;
		#400 //150996910000.0 * 2.7329482e+20 = 5.5250554e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111100000111100001100101101010;
		b = 32'b01010001000001100010011101001110;
		correct = 32'b01101010100101101101100011101101;
		#400 //3.2835934e+36 * 36011565000.0 = 9.118164e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111101110011011100001001100100;
		b = 32'b01101101001110110011111110111111;
		correct = 32'b11010000000011001010011101000000;
		#400 //-3.4187634e+37 * 3.6219226e+27 = -9439085000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010101011001010011110100110110;
		b = 32'b10011101010010110001010000011100;
		correct = 32'b00110111100100000111110100101011;
		#400 //-4.629447e-26 * -2.6877223e-21 = 1.7224424e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000101110001001101011110000001;
		b = 32'b11010001100010110000111110111110;
		correct = 32'b10110011101101010010111100101011;
		#400 //6298.938 * -74658070000.0 = -8.437049e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100100100110101101101011100100;
		b = 32'b00111110110110101100010101001010;
		correct = 32'b00100101001101010011010100100001;
		#400 //6.715767e-17 * 0.42728645 = 1.5717248e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001010000011001011000100010111;
		b = 32'b11101100011010001010010111000101;
		correct = 32'b10011101000110101101000001100001;
		#400 //2305093.8 * -1.12501446e+27 = -2.048946e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101010110000111100100100001011;
		b = 32'b01100101011011000000110011010110;
		correct = 32'b01000100110101000101010100001010;
		#400 //1.1834497e+26 * 6.9669704e+22 = 1698.6575
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110001001110011011000110111;
		b = 32'b10001010010000010001110011100111;
		correct = 32'b11110011010111011010101000001000;
		#400 //0.16329275 * -9.298048e-33 = -1.7562046e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101011010001101010011001101011;
		b = 32'b10011110110001111100100000101110;
		correct = 32'b01001011111111101000110010110011;
		#400 //-7.057468e-13 * -2.1152737e-20 = 33364326.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100101001000001111011100110100;
		b = 32'b00100110010010100011011011100000;
		correct = 32'b01111110010010111100011110100010;
		#400 //4.750867e+22 * 7.01572e-16 = 6.771746e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001100010000100010000011100010;
		b = 32'b00101001110111011000101100001001;
		correct = 32'b10100001111000000101001001001110;
		#400 //-1.4955112e-31 * 9.83849e-14 = -1.5200616e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010011111111010010111000101110;
		b = 32'b11001010110010011100110100111000;
		correct = 32'b01001000101000001001011010111110;
		#400 //-2174803000000.0 * -6612636.0 = 328885.94
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100001000001010110011110000010;
		b = 32'b11100101001101010000000100011111;
		correct = 32'b00111011001111001010110110000100;
		#400 //-1.5380472e+20 * -5.3423063e+22 = 0.0028789947
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111011001001100001000100010000;
		b = 32'b01101001100011111000010100110101;
		correct = 32'b00010001000101000001101110101111;
		#400 //0.002533976 * 2.168818e+25 = 1.1683672e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100101000010100000001011011000;
		b = 32'b00001100101111010101111010001000;
		correct = 32'b01010111101110101001001000111000;
		#400 //1.1970555e-16 * 2.9176955e-31 = 410274340000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110000000011101111010010110101;
		b = 32'b11010011011111100011100111001101;
		correct = 32'b01011100000011111111010000011101;
		#400 //-1.7697082e+29 * -1091891400000.0 = 1.620773e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111010000011010111001111111110;
		b = 32'b00010111101001010101010110001010;
		correct = 32'b01100001110110110000010111101001;
		#400 //0.00053960073 * 1.0684468e-24 = 5.0503285e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010111010110001110110011110011;
		b = 32'b10010111101101101110000010101010;
		correct = 32'b11111111000101111101010010111000;
		#400 //238512200000000.0 * -1.1818188e-24 = -2.0181793e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111010001010000001110101011001;
		b = 32'b11111001100010101010100010111011;
		correct = 32'b01000000000110110011000011110011;
		#400 //-2.1822528e+35 * -8.99949e+34 = 2.4248626
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111010101110010000100000010101;
		b = 32'b00011010100110111000110110101000;
		correct = 32'b01011111100110000100000110111000;
		#400 //0.0014116789 * 6.4335355e-23 = 2.1942505e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001010111110100010011100111111;
		b = 32'b10101010110111111000000100101000;
		correct = 32'b00011111100011110100001011111011;
		#400 //-2.4088887e-32 * -3.9702378e-13 = 6.0673666e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101000010101111000000010000101;
		b = 32'b01001101100001011001101101100010;
		correct = 32'b11011010010011100111010101010000;
		#400 //-4.0707182e+24 * 280194100.0 = -1.4528208e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001000110110000101011101000100;
		b = 32'b00100011000110000101110001010100;
		correct = 32'b11100101001101011100000000100100;
		#400 //-443066.12 * 8.259488e-18 = -5.3643294e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100010110111011101000101110110;
		b = 32'b00101100100010111111010111000010;
		correct = 32'b00110101110010101101110011111010;
		#400 //6.0123945e-18 * 3.977902e-12 = 1.5114485e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010011101101010000001001000101;
		b = 32'b00111100011001001011011111100101;
		correct = 32'b11010110110010101001100110000111;
		#400 //-1554854300000.0 * 0.0139598595 = -111380370000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000110101001001000010100110110;
		b = 32'b01001001010111001110110011110100;
		correct = 32'b00111100101111101010001111001010;
		#400 //21058.605 * 904911.25 = 0.02327146
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011010110111101111000100101000;
		b = 32'b00010000010100101100101000100010;
		correct = 32'b01001010000001110110000100100100;
		#400 //9.220666e-23 * 4.1570915e-29 = 2218057.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101111111101101000111111110100;
		b = 32'b00100001100001101100011100001010;
		correct = 32'b01001101111010100010100111011110;
		#400 //4.4849424e-10 * 9.132878e-19 = 491076540.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111000100110010110001010101101;
		b = 32'b11101101101011100011001010111010;
		correct = 32'b10001010011000010110100111110010;
		#400 //7.313988e-05 * -6.7389645e+27 = -1.0853282e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011100011110011000010100010101;
		b = 32'b00111110110011101111011010010100;
		correct = 32'b10011101000110100101000111100101;
		#400 //-8.2559194e-22 * 0.404225 = -2.0424069e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111011111110111111001010010100;
		b = 32'b10111001101111101000000100000110;
		correct = 32'b11000001101010010100100010111000;
		#400 //0.0076888297 * -0.00036335754 = -21.160507
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010001001000000101111001001000;
		b = 32'b00111010010110110010110001101000;
		correct = 32'b01010110001110110101000001101001;
		#400 //43048534000.0 * 0.0008360804 = 51488510000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011010110110001110100000101011;
		b = 32'b00000101000101110100101000010101;
		correct = 32'b11010101001101111000010000110011;
		#400 //-8.9710594e-23 * 7.1135926e-36 = -12611151000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001000100000001011101010101001;
		b = 32'b00100000011100010111010010000001;
		correct = 32'b01100111100010000111101111001101;
		#400 //263637.28 * 2.0452042e-19 = 1.2890511e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110100101110100110101101101;
		b = 32'b00111010011001110110110100010010;
		correct = 32'b01000011101001110101111001010100;
		#400 //0.2955126 * 0.00088282034 = 334.73694
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100100111101101001100011110011;
		b = 32'b01001110010101101111010010000001;
		correct = 32'b01010110000100101101011110011001;
		#400 //3.6391362e+22 * 901587000.0 = 40363670000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100001110000110001011101111001;
		b = 32'b10101001000101100101111101011001;
		correct = 32'b10111000001001100001000011011111;
		#400 //1.3219927e-18 * -3.338939e-14 = -3.9593197e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001001100001111011110100100111;
		b = 32'b00010100000010000110010011011101;
		correct = 32'b00110100111111101100010100111001;
		#400 //3.2677946e-33 * 6.886137e-27 = 4.7454685e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001001111001110001000100100010;
		b = 32'b01101111100001000000101101100101;
		correct = 32'b00011001110111111111110101000111;
		#400 //1892900.2 * 8.173159e+28 = 2.3159957e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001101111100101100011000000101;
		b = 32'b01011001001001101101111101110010;
		correct = 32'b00110100001110100011100000111111;
		#400 //509132960.0 * 2935658000000000.0 = 1.7343062e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010100111101101001011011001110;
		b = 32'b00110100101101111101000111100000;
		correct = 32'b10011111101010111011010101011000;
		#400 //-2.4899134e-26 * 3.423911e-07 = -7.2721325e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110110000001000001010000001000;
		b = 32'b11101110011110110110000100110110;
		correct = 32'b01000111000001101000000101111100;
		#400 //-6.697163e+32 * -1.9449565e+28 = 34433.484
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110010000001010100110101001111;
		b = 32'b10110101100100001111001100010010;
		correct = 32'b10111011111010110110110111010000;
		#400 //7.759197e-09 * -1.0799579e-06 = -0.0071847215
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100001001110110000100001000110;
		b = 32'b01000011001101101110110111100110;
		correct = 32'b01011101100000101101111011111001;
		#400 //2.1563358e+20 * 182.92929 = 1.178781e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001110111101000010011110111011;
		b = 32'b10010100010111001010100110110101;
		correct = 32'b11111010000011011010000010001110;
		#400 //2048122200.0 * -1.114063e-26 = -1.8384257e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001011011111010100101101111101;
		b = 32'b10011101111010000000000111111111;
		correct = 32'b11101101000010111011111010000100;
		#400 //16599933.0 * -6.1411953e-21 = -2.703046e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001011101100110100110000101111;
		b = 32'b10010000010101101011101000001010;
		correct = 32'b11111010110101011100001011001101;
		#400 //23500894.0 * -4.2347378e-29 = -5.5495513e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001011100110111110001011011110;
		b = 32'b01100011001011000101101110100011;
		correct = 32'b00100111111001111000100011101010;
		#400 //20432316.0 * 3.179443e+21 = 6.4263822e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001111001001010111011001100010;
		b = 32'b01001010100111001010101100100111;
		correct = 32'b00000100000001110010111101001000;
		#400 //8.157928e-30 * 5133715.5 = 1.5890884e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100101110011101110011000011010;
		b = 32'b01011001101010101100110100111100;
		correct = 32'b00001011100110110000110100101100;
		#400 //3.5891226e-16 * 6009550500000000.0 = 5.972365e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010000101001100000001001101000;
		b = 32'b00011001110111110001101000110111;
		correct = 32'b10110110001111100111110100000100;
		#400 //-6.547916e-29 * 2.3068248e-23 = -2.8384975e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000110011000001110100111000001;
		b = 32'b10111001001100010001000111110100;
		correct = 32'b11001100101000101001010110101001;
		#400 //14394.438 * -0.00016886723 = -85241160.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100011011111001000001000101010;
		b = 32'b00001001101100011101110101110010;
		correct = 32'b01011001001101011011011110000111;
		#400 //1.3688511e-17 * 4.2819446e-33 = 3196797600000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000100110011111101010110101101;
		b = 32'b10111000100110101101000110100001;
		correct = 32'b00001011101010111101010011111111;
		#400 //-4.8861696e-36 * -7.382339e-05 = 6.6187285e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010110010101000000110000100111;
		b = 32'b10111010001101101011001000110011;
		correct = 32'b11011011100101001001000001100111;
		#400 //58287165000000.0 * -0.0006969303 = -8.363414e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101101110000111010101101110000;
		b = 32'b10010011110111010100001011001000;
		correct = 32'b01011001011000100110010000001111;
		#400 //-2.2245067e-11 * -5.5854095e-27 = 3982710000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101010001011010000111011010110;
		b = 32'b11010001011011111011000001111010;
		correct = 32'b10011000001110001101010110011010;
		#400 //1.5370634e-13 * -64341123000.0 = -2.3889284e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111010000011001101011000101000;
		b = 32'b00100110010011011011100100010110;
		correct = 32'b01010011001011110100000101111111;
		#400 //0.0005372488 * 7.13745e-16 = 752718100000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001111110111111101100000001101;
		b = 32'b01011010011110100000100111110001;
		correct = 32'b00110100111001010010111000111100;
		#400 //7510956500.0 * 1.7594919e+16 = 4.2688214e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111000100010010011111011000111;
		b = 32'b00001001110101000000001011001000;
		correct = 32'b11101110001001011011100010111010;
		#400 //-6.544362e-05 * 5.103976e-33 = -1.2822087e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010000100110100000011110000110;
		b = 32'b10000101000011100100010000000010;
		correct = 32'b11001011000010101001010110001001;
		#400 //6.075388e-29 * -6.689299e-36 = -9082249.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100001000000110010011101101100;
		b = 32'b10010001100010001100000101011110;
		correct = 32'b11001110111101011000001110111000;
		#400 //4.44367e-19 * -2.1576188e-28 = -2059525100.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100010010010100001010110101110;
		b = 32'b00000110010111111000100101100001;
		correct = 32'b11011011011001110110111011000011;
		#400 //-2.7387582e-18 * 4.2042569e-35 = -6.5142503e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011011001011110001110101111;
		b = 32'b11100011001101010101101011100100;
		correct = 32'b00100111101000100100000101100100;
		#400 //-15066031.0 * -3.34541e+21 = 4.503493e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110010010010110111111100101000;
		b = 32'b11101100000000001100011000111000;
		correct = 32'b10000101110010100100010111101011;
		#400 //1.1845067e-08 * -6.227143e+26 = -1.9021673e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110101100110101100111101110011;
		b = 32'b11100111010010010110010011101101;
		correct = 32'b10001101110001001100100100010001;
		#400 //1.153427e-06 * -9.510574e+23 = -1.2127838e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010001001010101010110001011101;
		b = 32'b11010111010100110110010101110010;
		correct = 32'b00111001010011101010111101000101;
		#400 //-45814764000.0 * -232432660000000.0 = 0.00019710984
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000001001110110001100000011111;
		b = 32'b11011101111010000001001011100111;
		correct = 32'b00100010110011100110001000010100;
		#400 //-11.693389 * -2.0903353e+18 = 5.5940256e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010011000000001110111011011000;
		b = 32'b01110100110001010010100010010010;
		correct = 32'b10011101101001110110100110101010;
		#400 //-553762950000.0 * 1.2496403e+32 = -4.4313786e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010111101110011000000101000001;
		b = 32'b10101100100110001101001110001000;
		correct = 32'b11101010100110110101111010111011;
		#400 //407929600000000.0 * -4.3435845e-12 = -9.391543e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000100000010111001100110101101;
		b = 32'b00010100111000000001001011000001;
		correct = 32'b11101110100111110111110110110100;
		#400 //-558.4012 * 2.2625617e-26 = -2.468004e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011001010000101010101011110010;
		b = 32'b10110011011000011101000111001011;
		correct = 32'b10100101010111001010111101010011;
		#400 //1.0064087e-23 * -5.25777e-08 = -1.914136e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000100000011100110111100010100;
		b = 32'b10011010101111110011111001001101;
		correct = 32'b10101000101111101010100111001010;
		#400 //1.6743024e-36 * -7.90964e-23 = -2.1167872e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100001001110100001101100101011;
		b = 32'b00110010011111010100101010110111;
		correct = 32'b00101110001111000001100010001111;
		#400 //6.305521e-19 * 1.4743526e-08 = 4.2768063e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101110101110010100010101010111;
		b = 32'b01001100000010101001010001110010;
		correct = 32'b11100010001010110010000001011010;
		#400 //-2.8669277e+28 * 36327880.0 = -7.891811e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110011100111001111110000011110;
		b = 32'b01001001110010101100000110101000;
		correct = 32'b10101001010001100011010101110100;
		#400 //-7.310176e-08 * 1660981.0 = -4.4011195e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101011101001011010111101111011;
		b = 32'b10100111010110101001111110111101;
		correct = 32'b01000011110000100000001011011000;
		#400 //-1.1772661e-12 * -3.0340172e-15 = 388.02222
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001110011001010010101000000001;
		b = 32'b11011000101000000110001101101100;
		correct = 32'b10110101001101101110001100101001;
		#400 //961183800.0 * -1410791000000000.0 = -6.8130845e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011001011101001010111010110100;
		b = 32'b00111101000011000100001010010010;
		correct = 32'b01011011110111110100101101111111;
		#400 //4304499000000000.0 * 0.034243174 = 1.2570386e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111101011101100000011011101000;
		b = 32'b00101001001111110001011001011110;
		correct = 32'b01010011101001001100110100100100;
		#400 //0.06006518 * 4.242992e-14 = 1415632700000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100101111100111010011000010110;
		b = 32'b01101001011111100100101110001111;
		correct = 32'b10111011111101010100100001000001;
		#400 //-1.4382485e+23 * 1.9213998e+25 = -0.00748542
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010101111001000111101000101011;
		b = 32'b00110110000100000100000011010000;
		correct = 32'b00011111010010101011110000000011;
		#400 //9.2281214e-26 * 2.1495398e-06 = 4.2930683e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110001011011000000110100001111;
		b = 32'b10101000101101000110111001010110;
		correct = 32'b01001000001001110111010100100001;
		#400 //-3.4349943e-09 * -2.0031865e-14 = 171476.52
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101110000011111010000010001100;
		b = 32'b01011111110011100101110010110100;
		correct = 32'b11001101101100100010110011000101;
		#400 //-1.1112611e+28 * 2.9739916e+19 = -373659800.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000010101011011101100100000101;
		b = 32'b01011101110110010110100100011010;
		correct = 32'b00100100010011001011010001111001;
		#400 //86.92387 * 1.9582602e+18 = 4.4388315e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110001000100000101111111110011;
		b = 32'b01111011100111101101101110100010;
		correct = 32'b10110100111010001010100100001111;
		#400 //-7.149094e+29 * 1.6496752e+36 = -4.3336374e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000110000010100111000100011001;
		b = 32'b00011110100101000101100100111100;
		correct = 32'b10100110111011101110011101111010;
		#400 //-2.6038006e-35 * 1.5707016e-20 = -1.6577309e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110011000001111001001100011;
		b = 32'b10000111000010011110001111111111;
		correct = 32'b01101110110100001100111111010101;
		#400 //-3.3519689e-06 * -1.0373736e-34 = 3.2312068e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011101101001010001100101010000;
		b = 32'b11111000001001101111100000011011;
		correct = 32'b10100100111111010010000111101000;
		#400 //1.4870785e+18 * -1.3546148e+34 = -1.097787e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000000000001111011001011101101;
		b = 32'b00101101110010001111111110001110;
		correct = 32'b01010001101011001101010011111100;
		#400 //2.1202958 * 2.2850857e-11 = 92788460000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000100110001110001100010000101;
		b = 32'b11000101101101101000111011000111;
		correct = 32'b00111110100010111001100001111011;
		#400 //-1592.7662 * -5841.847 = 0.2726477
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101101101101011100000001011001;
		b = 32'b11111000010110001101011101111110;
		correct = 32'b00110100110101101001001010100100;
		#400 //-7.031165e+27 * -1.7592294e+34 = 3.99673e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010000101101101000011101000010;
		b = 32'b10111110000010011010111100011110;
		correct = 32'b01010010001010011011000010101110;
		#400 //-24498540000.0 * -0.13445708 = 182203420000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011001001000000000001000010000;
		b = 32'b10000101010010001010100000111010;
		correct = 32'b01010011010011000010001110111011;
		#400 //-8.272223e-24 * -9.434853e-36 = 876772800000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011000000010010101111011110000;
		b = 32'b11000010011111000110101101100100;
		correct = 32'b01010101000010110101000111000101;
		#400 //-604163400000000.0 * -63.104874 = 9573957000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100001101011001111001101111101;
		b = 32'b01111000111000101010011110001110;
		correct = 32'b00101000010000110101011111110000;
		#400 //3.9879815e+20 * 3.6776797e+34 = 1.0843743e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011101010101101110111001100010;
		b = 32'b10111110110010000011101111001010;
		correct = 32'b11011110000010010110010101000000;
		#400 //9.67964e+17 * -0.39108115 = -2.4750974e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111101010100001110001001101001;
		b = 32'b11001111000010100010001110100110;
		correct = 32'b11101101110000011000110101110100;
		#400 //1.7353438e+37 * -2317592000.0 = -7.4877017e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111001010110011110000001101111;
		b = 32'b11011001111000010110111110010010;
		correct = 32'b10011110111101110110101010000000;
		#400 //0.0002077834 * -7931818000000000.0 = -2.619619e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010101001000000110011000000111;
		b = 32'b00001100001101010011100001011010;
		correct = 32'b11001000011000101001011000100011;
		#400 //-3.2392228e-26 * 1.396069e-31 = -232024.55
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001111110001000110010001111100;
		b = 32'b10101011010000111110001011000111;
		correct = 32'b00100100000000000101010011000010;
		#400 //-1.9365797e-29 * -6.9592634e-13 = 2.7827368e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111100001110100000000011101110;
		b = 32'b11011101110001010001011010010001;
		correct = 32'b10011101111100011001101000101001;
		#400 //0.011352761 * -1.7752122e+18 = -6.3951567e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001000110001101000000101111100;
		b = 32'b10010110011110001011001111001011;
		correct = 32'b01110001110011000101010010100000;
		#400 //-406539.88 * -2.0090013e-25 = 2.0235919e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001011001100101111000001001001;
		b = 32'b10100011001001101111011010100100;
		correct = 32'b11100111100010010010111000111011;
		#400 //11726921.0 * -9.051106e-18 = -1.295634e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011110000001001001100000010101;
		b = 32'b01011100110010011111100101101010;
		correct = 32'b11000000101010000000111110111001;
		#400 //-2.3886024e+18 * 4.5480563e+17 = -5.2519193
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010110100001000100010010100001;
		b = 32'b11010010101000111001101111100001;
		correct = 32'b01000011010011101111010111110111;
		#400 //-72715150000000.0 * -351347440000.0 = 206.9608
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100101111100010000001010011010;
		b = 32'b11110010100101100010100011010011;
		correct = 32'b10110010110011010111000110001111;
		#400 //1.4226729e+23 * -5.9484294e+30 = -2.3916781e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110011100010010100010000111111;
		b = 32'b11010011110101010011111001110100;
		correct = 32'b10011111001001001100100111111000;
		#400 //6.3919735e-08 * -1831751600000.0 = -3.4895415e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010110011101010001000110110111;
		b = 32'b10101000110010111001010101111010;
		correct = 32'b00101101000110100001010101001101;
		#400 //-1.9796532e-25 * -2.2602353e-14 = 8.758616e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011000000001101011110110010101;
		b = 32'b11100100111100111000010010011110;
		correct = 32'b10110010100011011010010110011101;
		#400 //592595200000000.0 * -3.593692e+22 = -1.6489873e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100100011011011100111110100001;
		b = 32'b00011001001100000001111010111011;
		correct = 32'b11001010101011001101010111101010;
		#400 //-5.156705e-17 * 9.105193e-24 = -5663477.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100111111000101000111100111;
		b = 32'b11010110011010101110010011100100;
		correct = 32'b10101110000010010111111011101100;
		#400 //2018.5594 * -64567200000000.0 = -3.1262923e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000010000000110110000110011001;
		b = 32'b10011000101111101111000111010111;
		correct = 32'b00101000101100000010010010100101;
		#400 //-9.652369e-38 * -4.9358045e-24 = 1.9555817e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011101001101011110011110010111;
		b = 32'b01001101100111010010100010001000;
		correct = 32'b11001111000101000010011110101111;
		#400 //-8.192257e+17 * 329584900.0 = -2485628700.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111011010000011000110011000001;
		b = 32'b11101101001111001111011001010010;
		correct = 32'b10001101100000110001101110001011;
		#400 //0.0029533359 * -3.6550603e+27 = -8.080129e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111010111110110110110100010101;
		b = 32'b01111100100111000000111110100011;
		correct = 32'b10111101110011100011011110110100;
		#400 //-6.5273948e+35 * 6.4825237e+36 = -0.10069218
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100011010110000001001000100011;
		b = 32'b10111010010111010001010101010011;
		correct = 32'b11101000011110100011001000100111;
		#400 //3.9858036e+21 * -0.00084336585 = -4.726067e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110011001110010110010101011111;
		b = 32'b11001100101111011000001011101110;
		correct = 32'b01100101111110100111000011001111;
		#400 //-1.4688583e+31 * -99358580.0 = 1.4783407e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010010011001101010100001111010;
		b = 32'b00001100101000111100101001001000;
		correct = 32'b01000101001101000100000110101001;
		#400 //7.2782867e-28 * 2.523587e-31 = 2884.1038
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011001010110110011001011010111;
		b = 32'b11011110110100101101111100101101;
		correct = 32'b10111010000001010000110111101110;
		#400 //3856182400000000.0 * -7.5974566e+18 = -0.0005075623
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110010001011111010111000011;
		b = 32'b11100010110100011010011000100010;
		correct = 32'b10011010111100011011101000001101;
		#400 //0.19332032 * -1.9336703e+21 = -9.9975845e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101110000010111000101011111101;
		b = 32'b01100111110100101101110010101100;
		correct = 32'b10000101101010010110101000000000;
		#400 //-3.1728387e-11 * 1.9915353e+24 = -1.5931622e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011100011101100000110010001000;
		b = 32'b00111000101111110000010110100011;
		correct = 32'b01100011001001001101111101011000;
		#400 //2.7702649e+17 * 9.10864e-05 = 3.0413596e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011100010111011001110111100001;
		b = 32'b00100111000011000100001110111110;
		correct = 32'b11110100110010100011110100011110;
		#400 //-2.4951824e+17 * 1.9465626e-15 = -1.2818403e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000101111010010010111011010001;
		b = 32'b10000110101000100110010011110111;
		correct = 32'b11111110101101111100101110111010;
		#400 //7461.852 * -6.108598e-35 = -1.2215327e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001000100001010011100100101000;
		b = 32'b10110100101110000000011111011101;
		correct = 32'b10010011001110010101001010111011;
		#400 //8.018084e-34 * -3.4278392e-07 = -2.3391072e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011000101000000011101101110;
		b = 32'b00110100100101011100100100000001;
		correct = 32'b11010101111111001111111110100000;
		#400 //-9701230.0 * 2.7899662e-07 = -34771854000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010011000101010111000110000011;
		b = 32'b00111110011111010000101011011100;
		correct = 32'b00010100000101110011000010101011;
		#400 //1.886241e-27 * 0.24711174 = 7.63315e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110110011110110101100101101011;
		b = 32'b11000011110110111100001100010001;
		correct = 32'b11110010000100100110010111100010;
		#400 //1.2744923e+33 * -439.52396 = -2.8997107e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110001111001011100100000011010;
		b = 32'b11101011111111110011101001110110;
		correct = 32'b01000101011001100111100111110010;
		#400 //-2.2756472e+30 * -6.171043e+26 = 3687.6216
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001011001111100110110111110110;
		b = 32'b00110011011001110000001100110001;
		correct = 32'b01010111010100110000011100000100;
		#400 //12479990.0 * 5.378678e-08 = 232027090000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010101101110010000011101000110;
		b = 32'b01001010111111011001110000011100;
		correct = 32'b01001010001110101100010110110010;
		#400 //25430111000000.0 * 8310286.0 = 3060076.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101111000101101000110110011100;
		b = 32'b01010111011110010000010000110100;
		correct = 32'b11010111000110101100011001111111;
		#400 //-4.6593947e+28 * 273796450000000.0 = -170177320000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100111110000100110010010011000;
		b = 32'b11010011110000010000010011110000;
		correct = 32'b10010011100000001110100100110011;
		#400 //5.395488e-15 * -1658023000000.0 = -3.2541695e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001100000000111011111101000100;
		b = 32'b01000101011101111110010110010110;
		correct = 32'b01000110000010000000110110111100;
		#400 //34536720.0 * 3966.349 = 8707.434
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101010000110100101001010101001;
		b = 32'b00101100101010111000000011001111;
		correct = 32'b11111100111001100101101011110100;
		#400 //-4.664123e+25 * 4.874413e-12 = -9.568584e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000111011100001011000011000011;
		b = 32'b10110000001001010101111100111111;
		correct = 32'b10010110101110100100110000100001;
		#400 //1.8107539e-34 * -6.0162003e-10 = -3.0097965e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010000010000101011011010110110;
		b = 32'b00111010110010111000101001100000;
		correct = 32'b01010100111101001110010111110001;
		#400 //13067016000.0 * 0.001552891 = 8414638400000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110101100100111000011000111111;
		b = 32'b10100011111011111011000000011100;
		correct = 32'b11010001000111011001000001110010;
		#400 //1.0991424e-06 * -2.5987017e-17 = -42295830000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101001101010110000101001111011;
		b = 32'b10111001110010001101100101011110;
		correct = 32'b11101111010110100000000111000010;
		#400 //2.5846976e+25 * -0.00038308924 = -6.7469857e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000001110100000011101100110010;
		b = 32'b10000111101011111111110100010101;
		correct = 32'b01111001100101110111001101100001;
		#400 //-26.028904 * -2.6479822e-34 = 9.829712e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111001111110001011101011111011;
		b = 32'b01101110110010101101011010011001;
		correct = 32'b00001010100111001111010111000001;
		#400 //0.00047441557 * 3.1387702e+28 = 1.5114696e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010001111000000010110011000100;
		b = 32'b10010100011000110111001100011011;
		correct = 32'b10111100111111000101000001101110;
		#400 //3.5368558e-28 * -1.1483272e-26 = -0.03080007
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100100110101111101100001010000;
		b = 32'b11111001000111000100111111001011;
		correct = 32'b00101011001100001100000000011011;
		#400 //-3.1853095e+22 * -5.0726044e+34 = 6.279436e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111011000000010101011010000;
		b = 32'b10011001110011101110011110111011;
		correct = 32'b11101101000010101010110111010011;
		#400 //57386.812 * -2.1393496e-23 = -2.682442e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001011001010000010001101110010;
		b = 32'b10000110001000101101100001101110;
		correct = 32'b01000100100001000010100100010010;
		#400 //-3.238229e-32 * -3.062782e-35 = 1057.2834
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011010000001111000100101101011;
		b = 32'b00101100000100110010101101110001;
		correct = 32'b00101101011010111100001111000011;
		#400 //2.802835e-23 * 2.0914071e-12 = 1.3401671e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001111101011011100110000000011;
		b = 32'b01100111001100001001000010111011;
		correct = 32'b00100111111110111111110001110000;
		#400 //5831657000.0 * 8.338063e+23 = 6.994019e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100000001010111000000101100001;
		b = 32'b11000000111101100111110111011100;
		correct = 32'b11011110101100100001111100000101;
		#400 //4.943306e+19 * -7.7028637 = -6.4174915e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011110110011010100010010111001;
		b = 32'b11001010101110010100001101011010;
		correct = 32'b00010011100011011101001001100111;
		#400 //-2.1733642e-20 * -6070701.0 = 3.5800877e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010001100001011111000110010010;
		b = 32'b11000101111010100011100111001001;
		correct = 32'b10001011000100100110010100111001;
		#400 //2.113258e-28 * -7495.223 = -2.819473e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000010001010101111101111101100;
		b = 32'b00100010100101110111100111110100;
		correct = 32'b11011111000100000111101111111100;
		#400 //-42.746017 * 4.1057755e-18 = -1.0411192e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010000000001101100011111000111;
		b = 32'b11000101110011000101001100010011;
		correct = 32'b10001001101010001101111000010111;
		#400 //2.6580743e-29 * -6538.3843 = -4.065338e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011000010100010000010010101011;
		b = 32'b10111000101111001010000110100000;
		correct = 32'b11011111000011011101010101111111;
		#400 //919271900000000.0 * -8.9946436e-05 = -1.0220215e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101001101000011001001100010011;
		b = 32'b01100111111101011001111111001111;
		correct = 32'b11000001001010000110011001011001;
		#400 //-2.441645e+25 * 2.3198555e+24 = -10.524987
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011111100001110010011110001000;
		b = 32'b11101000011110110011111010011101;
		correct = 32'b10110110100010011011011001101001;
		#400 //1.9477805e+19 * -4.745876e+24 = -4.1041535e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100110111000011101001111000101;
		b = 32'b01100011001101110010110010001101;
		correct = 32'b10000011000111011100111000111011;
		#400 //-1.5669912e-15 * 3.3789644e+21 = -4.6374894e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000010101001111110111010101000;
		b = 32'b00111011000110000100100010010110;
		correct = 32'b00000111000011010010011101000000;
		#400 //2.4675427e-37 * 0.0023236624 = 1.0619196e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111111111010110010110001000011;
		b = 32'b10110010011100111110010100010000;
		correct = 32'b01111111111010110010110001000011;
		#400 //nan * -1.4196544e-08 = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010001010101010010110101101;
		b = 32'b11000001110000101000011111100010;
		correct = 32'b00110111111000001001000111001000;
		#400 //-0.0006509673 * -24.316349 = 2.6770766e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111111001110110011001001011001;
		b = 32'b01111000110110110011101111111110;
		correct = 32'b10000101110110101001011011110000;
		#400 //-0.731237 * 3.5572806e+34 = -2.0556067e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011000100111111110101001100000;
		b = 32'b10110111100000010100101101111000;
		correct = 32'b00100000100111100101000001101000;
		#400 //-4.1337195e-24 * -1.5413141e-05 = 2.681945e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111001011101010011001101010001;
		b = 32'b11101010101101101001010010010011;
		correct = 32'b11001110001010111110011010001000;
		#400 //7.9572097e+34 * -1.1036306e+26 = -721003000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110010001011101000010110011100;
		b = 32'b01110000100100100010100111011011;
		correct = 32'b01000001000110001101010110011001;
		#400 //3.4567626e+30 * 3.618833e+29 = 9.552148
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001111110001100000100111001100;
		b = 32'b11111000110111100101110101001101;
		correct = 32'b00010110011000111111111010000001;
		#400 //-6645061600.0 * -3.6080696e+34 = 1.8417221e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010011011010011011011011010010;
		b = 32'b11011100001111100000101110001011;
		correct = 32'b10110110100111010110100110000100;
		#400 //1003794600000.0 * -2.1397175e+17 = -4.6912483e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100101010011111001100101011011;
		b = 32'b00001001000100000010100101000110;
		correct = 32'b01011011101110000101001101111100;
		#400 //1.8006347e-16 * 1.7352776e-33 = 1.03766376e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100111111010101100101001101001;
		b = 32'b10101010010010100001111001011000;
		correct = 32'b10111101000101001011000011100101;
		#400 //6.51675e-15 * -1.7951732e-13 = -0.036301512
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011100011100000011101011100011;
		b = 32'b11110011011100010011001100100111;
		correct = 32'b00101000011111101111100010000000;
		#400 //-2.7047496e+17 * -1.9109818e+31 = 1.4153717e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010001110010011010010101100001;
		b = 32'b10010111101001000111010101111100;
		correct = 32'b01111001100111001111000101101101;
		#400 //-108257880000.0 * -1.0627909e-24 = 1.0186188e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010010101000111011110000101101;
		b = 32'b10011011101011011100110100011100;
		correct = 32'b01110110011100010010110001010000;
		#400 //-351618370000.0 * -2.8752998e-22 = 1.2228929e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000011001010000000110011111;
		b = 32'b01001101011111000011100101000010;
		correct = 32'b10100010011010000110111101100000;
		#400 //-8.331202e-10 * 264475680.0 = -3.1500824e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110101010101111010111001101000;
		b = 32'b01011001100010110000100000110000;
		correct = 32'b00011011010001101001000100111010;
		#400 //8.0347536e-07 * 4891753000000000.0 = 1.6425101e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100010111000101000000001001010;
		b = 32'b11010010000011001101010001001001;
		correct = 32'b10010000010011011101111000001100;
		#400 //6.1393254e-18 * -151214240000.0 = -4.060018e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110001000101111110110101110000;
		b = 32'b01000111111011111010101010010111;
		correct = 32'b10101000101000100100100000010110;
		#400 //-2.210836e-09 * 122709.18 = -1.8016875e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100111100010110101010011011011;
		b = 32'b11101000101100000000000010010011;
		correct = 32'b00111110010010101010100101001111;
		#400 //-1.3159485e+24 * -6.649177e+24 = 0.19791149
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100000101010110010110010111110;
		b = 32'b10110010000110100111110100001000;
		correct = 32'b00101110000011011101001101001010;
		#400 //-2.8998135e-19 * -8.992409e-09 = 3.224735e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010111100101010000101111111000;
		b = 32'b10110011001000010101101110110110;
		correct = 32'b00100011111011000111011110101001;
		#400 //-9.631921e-25 * -3.7569144e-08 = 2.563785e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100000111101011000001000000100;
		b = 32'b11110011110111011000111000111001;
		correct = 32'b10101100100011011101011010001010;
		#400 //1.4152565e+20 * -3.510688e+31 = -4.0312797e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000011011110010011010010011000;
		b = 32'b11101111001001100000011101011100;
		correct = 32'b00010011110000000010000000001001;
		#400 //-249.20544 * -5.138341e+28 = 4.8499203e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100000011011100000001111100111;
		b = 32'b11011101011101010001110111110110;
		correct = 32'b00000010011110001001010100111001;
		#400 //-2.0160675e-19 * -1.103909e+18 = 1.8262987e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101010100111000010010111111100;
		b = 32'b00011100111000110110110001101110;
		correct = 32'b11001101001011111100010011010110;
		#400 //-2.7737524e-13 * 1.5049628e-21 = -184307040.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010101110110110001000001011000;
		b = 32'b10001100010111101111100100111000;
		correct = 32'b01001000111110111000001011100001;
		#400 //-8.847918e-26 * -1.7177254e-31 = 515095.03
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110000111101000110001101011111;
		b = 32'b01100001000101111111000111000111;
		correct = 32'b00001111010011011110000000110101;
		#400 //1.778158e-09 * 1.7518002e+20 = 1.0150461e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010100101101001101001001001001;
		b = 32'b00111101100111010011010000100011;
		correct = 32'b11010110100100110011101011110101;
		#400 //-6212977000000.0 * 0.0767596 = -80940710000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001110100001100101100100110000;
		b = 32'b11110100100000111111110101110001;
		correct = 32'b10011001100000100100100101111111;
		#400 //1126996000.0 * -8.3658605e+31 = -1.347137e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010000001101001000000110101001;
		b = 32'b10110111000101101101101111100000;
		correct = 32'b11011000100110010010011110111110;
		#400 //12113585000.0 * -8.99189e-06 = -1347167800000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011000011011011001111001000100;
		b = 32'b00101010010100101110001101110111;
		correct = 32'b01101101100100000011100101000111;
		#400 //1045056000000000.0 * 1.8730665e-13 = 5.5793857e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011011011110111011000011110101;
		b = 32'b10111011101111100000010001110100;
		correct = 32'b01011111001010011000101101111110;
		#400 //-7.0844785e+16 * -0.0057988707 = 1.2216997e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011011111101111100011101110000;
		b = 32'b11111011011011010110001001011001;
		correct = 32'b00100000000001011001101011100011;
		#400 //-1.3948721e+17 * -1.2325691e+36 = 1.1316786e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110001101000001110100100110110;
		b = 32'b01000101010000101010001000001001;
		correct = 32'b01101011110100111010010101000111;
		#400 //1.5935852e+30 * 3114.1272 = 5.117277e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011111101000101011110110100000;
		b = 32'b01000001011001010111100011111100;
		correct = 32'b11011101101101011000110111000111;
		#400 //-2.345341e+19 * 14.342037 = -1.6352914e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111100001111011100100111110001;
		b = 32'b01111100101000010110101011011110;
		correct = 32'b10111111000101100111111101110000;
		#400 //-3.94176e+36 * 6.7050185e+36 = -0.58788204
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010011000011101101110100111001;
		b = 32'b10001010100010111000001101011100;
		correct = 32'b11001000000000110001001100010010;
		#400 //1.803199e-27 * -1.3434625e-32 = -134220.28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100011111011001111001111000;
		b = 32'b11101100000000000001001110110010;
		correct = 32'b10010111111111010111011101111000;
		#400 //1014.4761 * -6.1934205e+26 = -1.63799e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011010101111111110100111000011;
		b = 32'b00100100011100111001001111001111;
		correct = 32'b10110101110010011011001101101010;
		#400 //-7.937341e-23 * 5.2817424e-17 = -1.5027883e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111001001110001111010101111100;
		b = 32'b01101111001010100011010110011000;
		correct = 32'b00001001100010110001011110000111;
		#400 //0.00017639057 * 5.2677243e+28 = 3.3485158e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001000000000001110100111010011;
		b = 32'b00100001111100101100011000110101;
		correct = 32'b10100101100001111110111110101111;
		#400 //-3.879346e-34 * 1.6451023e-18 = -2.3581183e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110100011101000000101100011110;
		b = 32'b11110100101110010011001011100111;
		correct = 32'b00111111001010001010101110011110;
		#400 //-7.734045e+31 * -1.1738371e+32 = 0.6588687
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110011001011001111001100101111;
		b = 32'b11010101111010000110101100101010;
		correct = 32'b10011100101111100111111101100010;
		#400 //4.0268045e-08 * -31943370000000.0 = -1.2606073e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011100110010010001010101111111;
		b = 32'b00101100011001000101010101011011;
		correct = 32'b11101111111000010111001011100101;
		#400 //-4.5280084e+17 * 3.244813e-12 = -1.3954605e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010000100100001111001101100110;
		b = 32'b01101110000101000111111111101101;
		correct = 32'b00100001111110011110000111001000;
		#400 //19454964000.0 * 1.1489609e+28 = 1.693266e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011100011010010001100010110001;
		b = 32'b01110001011010111110111100111110;
		correct = 32'b10101010011111001110101110101001;
		#400 //-2.6244327e+17 * 1.16829125e+30 = -2.2463857e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001100111110001101100100110100;
		b = 32'b00100100101101101101000000010001;
		correct = 32'b11100111101011100011110001111000;
		#400 //-130468260.0 * 7.9282396e-17 = -1.6456144e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100011000001011001001001111000;
		b = 32'b11101111111011000110001011110010;
		correct = 32'b00110010100100001010011110101000;
		#400 //-2.4639711e+21 * -1.4631616e+29 = 1.6840048e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011001011100001101111111100101;
		b = 32'b11100011100101000110000000100001;
		correct = 32'b10110101010011111100101111111000;
		#400 //4237510600000000.0 * -5.47409e+21 = -7.741032e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010101110100111111110110001010;
		b = 32'b01001111100000000000011010100111;
		correct = 32'b11000101110100111111001010000110;
		#400 //-29135737000000.0 * 4295839000.0 = -6782.3154
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100101111111101101000011111111;
		b = 32'b00110100101101110011100100101111;
		correct = 32'b11110000101100100000001111010011;
		#400 //-1.5041705e+23 * 3.4128013e-07 = -4.4074364e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000000011110111100101110111110;
		b = 32'b10101001001010010100001110101001;
		correct = 32'b10010110101110110011101101110111;
		#400 //1.1368855e-38 * -3.7584224e-14 = -3.0249007e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100111111111110101000011010000;
		b = 32'b11001001110010011011111011011011;
		correct = 32'b11011101101000011111110011111110;
		#400 //2.4113884e+24 * -1652699.4 = -1.4590605e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010111100110111110110001001011;
		b = 32'b10111000110100001101000101101010;
		correct = 32'b00011110001111110010011101001011;
		#400 //-1.0076289e-24 * -9.957219e-05 = 1.0119581e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101100000111100110000011111100;
		b = 32'b00101011000101000100001011001100;
		correct = 32'b01000000100010001011110000111000;
		#400 //2.2506988e-12 * 5.267286e-13 = 4.272976
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111011000100000000001000001001;
		b = 32'b11010000010100010010001010000101;
		correct = 32'b00101010001100000100011101011110;
		#400 //-0.002197387 * -14034802000.0 = 1.56567e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010111110010111010110000111111;
		b = 32'b10101101000001101000110111011101;
		correct = 32'b01101010010000011100000001111101;
		#400 //-447881300000000.0 * -7.648518e-12 = 5.855792e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001010101010100000001011001010;
		b = 32'b10100110000001001110111011100111;
		correct = 32'b10100100001000111011001110100011;
		#400 //1.6371454e-32 * -4.6120473e-16 = -3.549715e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010001101110101111110101101001;
		b = 32'b01001000000101011100101001100111;
		correct = 32'b01001001000111111100100110101001;
		#400 //100389430000.0 * 153385.61 = 654490.56
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010011100000010000111000111000;
		b = 32'b00110110111111100010110001001000;
		correct = 32'b10011100000000011111101110110100;
		#400 //-3.25782e-27 * 7.574945e-06 = -4.300784e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101100001100011111111111110000;
		b = 32'b10110100011101010010010011011100;
		correct = 32'b11110111001110011110000111100001;
		#400 //8.60754e+26 * -2.2830812e-07 = -3.7701417e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001100110000110010011010111101;
		b = 32'b11010000010001010100000100000000;
		correct = 32'b10111011111111010100010101101111;
		#400 //102315496.0 * -13237486000.0 = -0.0077292244
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000010010001101111000110001111;
		b = 32'b01010111111100001001100101100011;
		correct = 32'b10101001110100111010110110010100;
		#400 //-49.735897 * 529083160000000.0 = -9.400393e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010000100000110111000101111001;
		b = 32'b11001110100111011010101011111100;
		correct = 32'b10000001010101010110101110000000;
		#400 //5.184522e-29 * -1322614300.0 = -3.919905e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010110101011010110011001011100;
		b = 32'b00010010010011111111001001111100;
		correct = 32'b01000011110101010111100000101001;
		#400 //2.8014255e-25 * 6.561657e-28 = 426.93875
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100011101101100010110000101111;
		b = 32'b01110001111100000110100110111111;
		correct = 32'b10110001010000011111101111001011;
		#400 //-6.7209824e+21 * 2.3809357e+30 = -2.8228324e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000000100100111100011011111101;
		b = 32'b10010101110010111000100000101000;
		correct = 32'b11101010001110011101111101100000;
		#400 //4.6180406 * -8.2205864e-26 = -5.6176534e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000101101001001000111111000000;
		b = 32'b00101101011010000000101101111111;
		correct = 32'b01010111101101011000110011001100;
		#400 //5265.9688 * 1.3190226e-11 = 399232650000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100011001100111101000111011001;
		b = 32'b11110110100011111000101001101100;
		correct = 32'b00101100001000000101100111101000;
		#400 //-3.3170883e+21 * -1.4556757e+33 = 2.2787276e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101101110001011010011000101011;
		b = 32'b00110101001000100110111110110101;
		correct = 32'b10111000000110111011111101100111;
		#400 //-2.24701e-11 * 6.051226e-07 = -3.7133137e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000011000110111100111000111100;
		b = 32'b00111010001010011111101000110001;
		correct = 32'b00001000011010101010011111111111;
		#400 //4.578715e-37 * 0.000648412 = 7.061429e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101111010011001110010010110101;
		b = 32'b01000111111100000010111110000100;
		correct = 32'b01100110110110100110001001010001;
		#400 //6.341143e+28 * 122975.03 = 5.1564476e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101000100101101001011000010100;
		b = 32'b00000100101100101111001100010100;
		correct = 32'b11100011010101110110110010100000;
		#400 //-1.6718431e-14 * 4.207083e-36 = -3.9738772e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001100100011101101111101111110;
		b = 32'b01011001111000011101000111111011;
		correct = 32'b00110010001000011111011110100000;
		#400 //74906610.0 * 7945343000000000.0 = 9.427737e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101100101001101111000000100100;
		b = 32'b10011000001000000011101010001111;
		correct = 32'b11010100000001010101110000011011;
		#400 //4.7446647e-12 * -2.070908e-24 = -2291103700000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111101111101110111000010001101;
		b = 32'b11100110010101100101100010010011;
		correct = 32'b01010111000100111100001100101100;
		#400 //-4.1112964e+37 * -2.5305508e+23 = 162466470000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000111110110011110010101111110;
		b = 32'b10000101010000111000001101110100;
		correct = 32'b11000010000011101010011101100001;
		#400 //3.2785414e-34 * -9.193e-36 = -35.663456
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111101010010100110111011001011;
		b = 32'b01110000000110001011111000111010;
		correct = 32'b00001100101010011010001111110001;
		#400 //0.049422067 * 1.8908677e+29 = 2.6137241e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101001110000001111000110111100;
		b = 32'b10011110110111111000100010010101;
		correct = 32'b01001010010111001111011111001001;
		#400 //-8.568447e-14 * -2.3667532e-20 = 3620338.2
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110001110011001101000010110000;
		b = 32'b10110111000000010011100110110000;
		correct = 32'b00111010010010101101111110000010;
		#400 //-5.9609064e-09 * -7.702431e-06 = 0.0007738994
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110000010111110100100110100100;
		b = 32'b11101100001001001000100010011011;
		correct = 32'b01000011101011011011010101000110;
		#400 //-2.7641673e+29 * -7.9563574e+26 = 347.4162
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101101110001001110011111011110;
		b = 32'b10111110001101001111001101000001;
		correct = 32'b11101111000010110100100101011100;
		#400 //7.6174215e+27 * -0.17670919 = -4.3107102e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111010101110000000001110010010;
		b = 32'b11100010100111010001111010101001;
		correct = 32'b01010111100101011110100011100101;
		#400 //-4.777275e+35 * -1.449174e+21 = 329655000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101111100010100100100010000001;
		b = 32'b11001001001111011101110110110010;
		correct = 32'b11100101101110100111001100101111;
		#400 //8.559317e+28 * -777691.1 = -1.1006062e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101010101010011110001101110000;
		b = 32'b01001010001100011110101100100110;
		correct = 32'b01011111111101000111001000011110;
		#400 //1.0269125e+26 * 2915017.5 = 3.5228348e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000000011010110110110011010000;
		b = 32'b10000011101101111010111111110011;
		correct = 32'b11111100001001000000110110000001;
		#400 //3.6785164 * -1.0796169e-36 = -3.4072423e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001010100110000100010100011100;
		b = 32'b00011000100010100000011101100110;
		correct = 32'b00110001100011010011010011010010;
		#400 //1.4663064e-32 * 3.5679634e-24 = 4.109645e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101100111010000011101110101110;
		b = 32'b10001000000001111000101001100111;
		correct = 32'b11100100010110110101000000101001;
		#400 //6.6004624e-12 * -4.0787776e-34 = -1.6182452e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110000001010001011101011000;
		b = 32'b11000110100011101110000110110110;
		correct = 32'b10110110111011100111010101011101;
		#400 //0.12997186 * -18288.855 = -7.1066156e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101011011111000101001101111111;
		b = 32'b11001001110000011001011111001000;
		correct = 32'b01100001001001101101010101010101;
		#400 //-3.050436e+26 * -1585913.0 = 1.9234573e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000101110100100001010101001111;
		b = 32'b10000000111000101110001011000100;
		correct = 32'b01000100011011010000101010010011;
		#400 //-1.9756133e-35 * -2.083617e-38 = 948.1652
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011111100001000000010011000001;
		b = 32'b01001101011001010000100111111110;
		correct = 32'b10010001100100111000111100010110;
		#400 //-5.591204e-20 * 240164830.0 = -2.3280694e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111100110110001110000111000011;
		b = 32'b10001000001111100111101110000011;
		correct = 32'b11110100000100011011110101100101;
		#400 //0.02647484 * -5.7321233e-34 = -4.6186793e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111100001111111101110011011010;
		b = 32'b01000010101111100110111110111011;
		correct = 32'b10111001000000001111010101101010;
		#400 //-0.01171037 * 95.21822 = -0.00012298455
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001101000001110101111010001011;
		b = 32'b01111100000001010001100011000000;
		correct = 32'b10010000100000100010111110000100;
		#400 //-141945010.0 * 2.76431e+36 = -5.134917e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010101100000101101110010110001;
		b = 32'b11011110010100100001011001101010;
		correct = 32'b00110110100111110111010111101011;
		#400 //-17985547000000.0 * -3.784601e+18 = 4.7522967e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010101110000011100111001001010;
		b = 32'b10101001011001100000000000111010;
		correct = 32'b00101011110101111011011010100110;
		#400 //-7.8277546e-26 * -5.1070456e-14 = 1.5327364e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101110110011101001010110011001;
		b = 32'b11000110010000001101110100100010;
		correct = 32'b10101000000010010001101100101000;
		#400 //9.394369e-11 * -12343.283 = -7.610916e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111011001110011111011101010;
		b = 32'b01001001011100000001010101111010;
		correct = 32'b10101101011101101001001101110001;
		#400 //-1.3783321e-05 * 983383.6 = -1.401622e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100000111001000100110000101100;
		b = 32'b00011110110100101001000111101110;
		correct = 32'b11000001100010101100011010101110;
		#400 //-3.867511e-19 * 2.229497e-20 = -17.347012
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100000011100000111101101111111;
		b = 32'b11011000000111011101110111111111;
		correct = 32'b00000111110000101111110000110000;
		#400 //-2.0369652e-19 * -694307170000000.0 = 2.9338098e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110000101011101001011101010110;
		b = 32'b10110110110001111011000101001101;
		correct = 32'b01111001010111111101001000011010;
		#400 //-4.3226677e+29 * -5.9513027e-06 = 7.2633973e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001111011101110100110110100111;
		b = 32'b01010000100000001100101001110100;
		correct = 32'b10111110011101011100100011100111;
		#400 //-4149061400.0 * 17286013000.0 = -0.2400242
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101001111100011100000111111101;
		b = 32'b11111001100001101100011001010110;
		correct = 32'b10101111111001011001101011110100;
		#400 //3.65334e+25 * -8.747381e+34 = -4.1764958e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110001010111111011101001111000;
		b = 32'b00000001101001001000010101100010;
		correct = 32'b11101111001011100001000001110101;
		#400 //-3.2556766e-09 * 6.043548e-38 = -5.3870287e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100111001000011010111001010011;
		b = 32'b00001101000110100110110010010111;
		correct = 32'b11011001100001100000001111011001;
		#400 //-2.243774e-15 * 4.7585624e-31 = -4715234700000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000110001010010000111101101101;
		b = 32'b00111101110101000010111011001111;
		correct = 32'b00000111110010111111100011101001;
		#400 //3.17967e-35 * 0.103604905 = 3.0690341e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000111101010011100011100101;
		b = 32'b10001001011011000100110000011111;
		correct = 32'b01100111000001001101010110100100;
		#400 //-1.7842267e-09 * -2.8443259e-33 = 6.2729335e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100111001001111010011011001001;
		b = 32'b10101010110110111011000010111001;
		correct = 32'b11111011110000110101110001000010;
		#400 //7.9171185e+23 * -3.902484e-13 = -2.0287382e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111011011100110011101101010101;
		b = 32'b01011101010001010100100101000011;
		correct = 32'b10011101100111011100111101000110;
		#400 //-0.0037114222 * 8.8849796e+17 = -4.177187e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010101100010000111110010010110;
		b = 32'b10011001111000011101011111100000;
		correct = 32'b10111011000110101011011000101111;
		#400 //5.5126525e-26 * -2.3351646e-23 = -0.0023607125
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100100111010000001101000100011;
		b = 32'b00011001101011101001110010001010;
		correct = 32'b11001010101010100010010011010011;
		#400 //-1.0065824e-16 * 1.8054404e-23 = -5575273.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011011110111001100110011001001;
		b = 32'b10111000011111101111001000100111;
		correct = 32'b00100010110111011011011001111110;
		#400 //-3.6528286e-22 * -6.078384e-05 = 6.009539e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110001010100101000010110101010;
		b = 32'b10111111111000110010010011000011;
		correct = 32'b01110000111011010100010001010101;
		#400 //-1.0424551e+30 * -1.7745594 = 5.8744445e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000011101010010110101110101110;
		b = 32'b00101110011011100000010110110100;
		correct = 32'b10010100101101100011011110000110;
		#400 //-9.957649e-37 * 5.412e-11 = -1.8399204e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011100001101101010111111011;
		b = 32'b00011000111000111110001001111110;
		correct = 32'b11110010000101110111100010100010;
		#400 //-17673206.0 * 5.8906823e-24 = -3.0001966e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111111000010000101101111010000;
		b = 32'b11001111000111101101001101100111;
		correct = 32'b00101111010110111100100101101100;
		#400 //-0.53265095 * -2664654600.0 = 1.9989493e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100110001011101101111010101000;
		b = 32'b11011101000000100101101111110111;
		correct = 32'b10001000101010111011010001111000;
		#400 //6.067013e-16 * -5.870858e+17 = -1.0334116e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010111110111111001100011001001;
		b = 32'b01001001110011001000010101101001;
		correct = 32'b00001101100010111111000001000101;
		#400 //1.4449606e-24 * 1675437.1 = 8.624379e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101001011100001000111000001111;
		b = 32'b00010011011001010001000100001000;
		correct = 32'b11010101100001100110101101101010;
		#400 //-5.341392e-14 * 2.891226e-27 = -18474487000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011101111101011000011111011011;
		b = 32'b01010111110110110111110011001010;
		correct = 32'b01000101100011110011000000010100;
		#400 //2.2115438e+18 * 482658020000000.0 = 4582.01
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011001100101010001111101101100;
		b = 32'b01010110101001101000110100001000;
		correct = 32'b11000010011001010011011000110100;
		#400 //-5246790000000000.0 * 91562330000000.0 = -57.302933
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110011010001110010100111111010;
		b = 32'b11001100110010101111000000111010;
		correct = 32'b01100101111110110011110100011100;
		#400 //-1.5779395e+31 * -106398160.0 = 1.4830516e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000011100101001000111000101010;
		b = 32'b00101010101011010110100001101010;
		correct = 32'b10011000010110110100111101111100;
		#400 //-8.7312975e-37 * 3.0803425e-13 = -2.8345216e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110111010011101010000001011111;
		b = 32'b00011001110000110010000101000010;
		correct = 32'b01011101000001111000101010011011;
		#400 //1.2315896e-05 * 2.017596e-23 = 6.104243e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000100110000001010110101001000;
		b = 32'b00000100011000111111110010011010;
		correct = 32'b00111111110110000101100111111111;
		#400 //4.5298117e-36 * 2.679971e-36 = 1.6902465
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000001010111011011100000001001;
		b = 32'b00100011010110110101101010000100;
		correct = 32'b00011101100000010110000101010111;
		#400 //4.0723328e-38 * 1.1891181e-17 = 3.4246663e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110010110000000100000100001011;
		b = 32'b10101011011001001010001011110100;
		correct = 32'b01000110110101110100001101100100;
		#400 //-2.238132e-08 * -8.1228015e-13 = 27553.695
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100101101000001000010111011110;
		b = 32'b10111100101111110101101111001000;
		correct = 32'b10101000010101101011111110000000;
		#400 //2.7846288e-16 * -0.023359194 = -1.1920911e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101010100110011100110010000000;
		b = 32'b11100000110000000000111011111010;
		correct = 32'b11001001010011010000000010101101;
		#400 //9.296569e+25 * -1.1071419e+20 = -839690.8
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101100101110001011010000011111;
		b = 32'b01100001011000000010001111010011;
		correct = 32'b01001010110100101111010101000010;
		#400 //1.7863436e+27 * 2.5841575e+20 = 6912673.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010101101111001011010000110001;
		b = 32'b00011011000110100111001111100110;
		correct = 32'b11111010000111000110001010010010;
		#400 //-25935263000000.0 * 1.277603e-22 = -2.0299939e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101000000001001100010101101100;
		b = 32'b00001111001010001100000110010011;
		correct = 32'b01011000010010010110100101010101;
		#400 //7.370281e-15 * 8.3203205e-30 = 885816940000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000011010011100001101101001111;
		b = 32'b01101101110100011000001101001010;
		correct = 32'b00010100111110111101011010001011;
		#400 //206.10667 * 8.105136e+27 = 2.5429145e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011010010001100111001111000000;
		b = 32'b01000010010110011110011000010010;
		correct = 32'b11010111011010010010011100101110;
		#400 //-1.3964828e+16 * 54.474678 = -256354480000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100101111100000000110000100111;
		b = 32'b01101001001101101000010010011110;
		correct = 32'b10111100001010000101100001101110;
		#400 //-1.4169902e+23 * 1.3790673e+25 = -0.0102749895
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111101011000011111111010100100;
		b = 32'b11101101101110011001111111000111;
		correct = 32'b10001111000110111101011010010001;
		#400 //0.055174485 * -7.180986e+27 = -7.683414e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000101100101101101111001011110;
		b = 32'b10010001110001101010101011010100;
		correct = 32'b11110011010000100110100001000011;
		#400 //4827.796 * -3.1344173e-28 = -1.5402531e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000001010101000110101011011001;
		b = 32'b10110111000010100110000101010010;
		correct = 32'b01001001110001000111101111001010;
		#400 //-13.276086 * -8.2481e-06 = 1609593.2
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011011101011110110011110100010;
		b = 32'b10111010010111011011111111110100;
		correct = 32'b00100000110010100111111100110000;
		#400 //-2.9018293e-22 * -0.0008459084 = 3.4304297e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001101101111101001001101001011;
		b = 32'b11101001010110100101111011011000;
		correct = 32'b00100011110111110110101001001101;
		#400 //-399665500.0 * -1.6499607e+25 = 2.4222729e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011010100000000001010111001010;
		b = 32'b11101001110010001010111110010111;
		correct = 32'b00110000001000110110001101111100;
		#400 //-1.8026377e+16 * -3.0326795e+25 = 5.944043e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100110110010001110100101011111;
		b = 32'b01010011101010101101110111110110;
		correct = 32'b01010010100101101000000111001011;
		#400 //4.743891e+23 * 1467736700000.0 = 323211330000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100111000000001011011111000011;
		b = 32'b10101010001100001000101011101100;
		correct = 32'b00111100001110101010011010000010;
		#400 //-1.7863186e-15 * -1.5680138e-13 = 0.011392238
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100110110001010110100100011110;
		b = 32'b01011010010100101010100111001110;
		correct = 32'b10001011111011111110010100101101;
		#400 //-1.3698113e-15 * 1.4824112e+16 = -9.2404277e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000110011001100011100000110010;
		b = 32'b11000001001101110000101101011111;
		correct = 32'b00000100101000001111110100100001;
		#400 //-4.3299478e-35 * -11.440276 = 3.784828e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010001001101000011011111110;
		b = 32'b00111000000111111111011101100001;
		correct = 32'b11000001100001010011111111111001;
		#400 //-0.0006352513 * 3.8138944e-05 = -16.656237
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101110000010110101010000010010;
		b = 32'b11011011000010101000101100111000;
		correct = 32'b00010010100000001011100110010001;
		#400 //-3.167961e-11 * -3.899662e+16 = 8.123681e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111010011101001010100111010011;
		b = 32'b11000010101111001110100101110011;
		correct = 32'b01110111001001011100011001110100;
		#400 //-3.1759122e+35 * -94.455956 = 3.3623207e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111100100011010000110010011000;
		b = 32'b01000010111101001010101111101111;
		correct = 32'b11111001000100111001010001101111;
		#400 //-5.858954e+36 * 122.33581 = -4.789239e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001111110101111000101001101100;
		b = 32'b11010010100010101100000100001001;
		correct = 32'b10111100110001101101010111011010;
		#400 //7232346000.0 * -297972040000.0 = -0.024271894
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010110011010001110011101011110;
		b = 32'b00100010101111010110010010010111;
		correct = 32'b01110011000111010110100000010010;
		#400 //64020103000000.0 * 5.1335056e-18 = 1.247103e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010011001100110101010010100011;
		b = 32'b01100111011010010111100010111000;
		correct = 32'b00101011010001001010001010000011;
		#400 //770219100000.0 * 1.10253826e+24 = 6.985872e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110001010101011101100101110100;
		b = 32'b00010011010100110010000000001101;
		correct = 32'b11011101100000011010011011010001;
		#400 //-3.1119187e-09 * 2.6647746e-27 = -1.167798e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111100110101101110100011010000;
		b = 32'b00010000111101010111000001010110;
		correct = 32'b11101011011000000010100000101101;
		#400 //-0.02623406 * 9.680854e-29 = -2.709891e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110011110010100100010101100010;
		b = 32'b10010001000001110001100000011110;
		correct = 32'b01100010001111111010011000101111;
		#400 //-9.418979e-08 * -1.0657054e-28 = 8.838257e+20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001111111100000011001001000110;
		b = 32'b01111001010111111111001010011001;
		correct = 32'b10010110000010010100100110000011;
		#400 //-8059653000.0 * 7.2675167e+34 = -1.1089968e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011000111011110000001000110001;
		b = 32'b00111101001101011010100010011010;
		correct = 32'b00011011001010000110100011101011;
		#400 //6.1782265e-24 * 0.044350244 = 1.3930535e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100010001011100111000100000010;
		b = 32'b11110101001101011110110100000011;
		correct = 32'b10101100011101010111011111011101;
		#400 //8.044691e+20 * -2.3061838e+32 = -3.4883132e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000011111000101111101011001101;
		b = 32'b11110011100010101111001001001000;
		correct = 32'b10001111110100010001100100001111;
		#400 //453.95938 * -2.2016938e+31 = -2.0618643e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100010001110000111111000101010;
		b = 32'b01010010110110001011111001011111;
		correct = 32'b00001110110110011110100001110000;
		#400 //2.500344e-18 * 465453420000.0 = 5.371846e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001101011110100110001011011001;
		b = 32'b10100011100011110100011010111111;
		correct = 32'b00101001010111111011000010000111;
		#400 //-7.715618e-31 * -1.5534053e-17 = 4.966906e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001010110101001001101000110110;
		b = 32'b00001111100000010111010001110001;
		correct = 32'b11111010110100100011011010001110;
		#400 //-6966555.0 * 1.2765234e-29 = -5.4574442e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100000001101010111011111110111;
		b = 32'b11110000001000000110110001010001;
		correct = 32'b10101111100100001100101011000000;
		#400 //5.2304766e+19 * -1.985942e+29 = -2.633751e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011100101101101001111101100110;
		b = 32'b00111000111000100010110001010001;
		correct = 32'b10100011010011101011010011001110;
		#400 //-1.2084953e-21 * 0.00010784774 = -1.1205569e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000000100111000011110111010111;
		b = 32'b10011010110101011110001100011111;
		correct = 32'b11100101001110110000000100011110;
		#400 //4.882549 * -8.846167e-23 = -5.5193946e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111100100010011001011101000011;
		b = 32'b10010110010010110111100101010001;
		correct = 32'b11100101101011010001110000001000;
		#400 //0.01679576 * -1.643649e-25 = -1.0218581e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100110011101101111001010111011;
		b = 32'b00010101011001111000110001110111;
		correct = 32'b11010000100010001000001101001000;
		#400 //-8.5677356e-16 * 4.6760886e-26 = -18322440000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101001101100111110110001111000;
		b = 32'b01010101011011111000010101111011;
		correct = 32'b00010011110000000100110101010110;
		#400 //7.9902176e-14 * 16459786000000.0 = 4.8543873e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100000111100000101100110010110;
		b = 32'b11101111011001010111000010010101;
		correct = 32'b10110001000001100001011000101010;
		#400 //1.3855231e+20 * -7.100817e+28 = -1.9512165e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100000111110101001101110101111;
		b = 32'b01100100110001101101111010110001;
		correct = 32'b10111011101000010100110011110111;
		#400 //-1.4446576e+20 * 2.9348015e+22 = -0.004922505
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101000000101110101000001010000;
		b = 32'b11001001000100100011110111000001;
		correct = 32'b10011110100001000111000010010110;
		#400 //8.399599e-15 * -599004.06 = -1.4022608e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010111111001110111011110110100;
		b = 32'b10101101110011110001000101011101;
		correct = 32'b01101001100011110001010100110101;
		#400 //-509002600000000.0 * -2.3540886e-11 = 2.1622067e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011101011000101110011110110001;
		b = 32'b10101101010111010011101000000100;
		correct = 32'b10101111100000110100100100010110;
		#400 //3.0030633e-21 * -1.2575278e-11 = -2.3880692e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011100010011110000110000101000;
		b = 32'b11111000001000110110001011011000;
		correct = 32'b10100011101000100011010010001001;
		#400 //2.3311474e+17 * -1.3255456e+34 = -1.7586325e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011101001111110010000010101001;
		b = 32'b00100001101001010101101000101000;
		correct = 32'b00111011000100111111001111110000;
		#400 //2.5295524e-21 * 1.1204699e-18 = 0.0022575818
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110011001010101111011110111110;
		b = 32'b00100100000011110001010011001011;
		correct = 32'b01001110100110001111001001111011;
		#400 //3.980653e-08 * 3.1025794e-17 = 1283014000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100100100001011000010010100110;
		b = 32'b00011011110001111010110011011110;
		correct = 32'b01001000001010110010111001100010;
		#400 //5.790427e-17 * 3.30335e-22 = 175289.53
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001001010110010011000111001000;
		b = 32'b01100101000001100101000110100001;
		correct = 32'b00100011110011101111101000010001;
		#400 //889628.5 * 3.964393e+22 = 2.2440472e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100010100011110100101110110101;
		b = 32'b10110101111000110111010001110001;
		correct = 32'b00101100001000010100011101110001;
		#400 //-3.8840386e-18 * -1.6946707e-06 = 2.2919134e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010100101001110000010111000110;
		b = 32'b11001010100011110000010110010011;
		correct = 32'b00001001100101010111101011011110;
		#400 //-1.6864968e-26 * -4686537.5 = 3.598599e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011100111110001011110100111101;
		b = 32'b11010001101010110010101011000100;
		correct = 32'b11001010101110100000001001010000;
		#400 //5.601109e+17 * -91894610000.0 = -6095144.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100011101010011011010011100111;
		b = 32'b00101100100111101011000011101111;
		correct = 32'b11110110100010001110001010010101;
		#400 //-6.26107e+21 * 4.5102737e-12 = -1.3881797e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110111101100100101111101000100;
		b = 32'b10011010001010100110000110000101;
		correct = 32'b11011101000001100000000011100010;
		#400 //2.1263615e-05 * -3.5233952e-23 = -6.034979e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100100010000100010001010011110;
		b = 32'b00111100101111001011010111010111;
		correct = 32'b10100111000000111010110111111110;
		#400 //-4.2096366e-17 * 0.023035927 = -1.8274223e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101000100010110101010001101011;
		b = 32'b00111011111010101111110111111011;
		correct = 32'b00101100000101111100100100011101;
		#400 //1.546871e-14 * 0.00717139 = 2.157003e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010100100111101111011001111000;
		b = 32'b00000100111010111001101000001000;
		correct = 32'b01001111001011001011100111001000;
		#400 //1.6051138e-26 * 5.538969e-36 = 2897856500.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010111001110011101100001010100;
		b = 32'b11001101100011100000111111101001;
		correct = 32'b10001001001001110111001011110001;
		#400 //6.004977e-25 * -297925920.0 = -2.0155939e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110110111001111000110011100101;
		b = 32'b01000001010011011011001000100000;
		correct = 32'b01110101000100000001011010110111;
		#400 //2.3481997e+33 * 12.855988 = 1.8265416e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010100010001000110110000010001;
		b = 32'b11011001101010101010100111001011;
		correct = 32'b10111010000100110101000111001110;
		#400 //3374506600000.0 * -6004679400000000.0 = -0.0005619795
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001010100100000110010011011110;
		b = 32'b00100110000111000011101010100001;
		correct = 32'b11100011111011001001101101011111;
		#400 //-4731503.0 * 5.420283e-16 = -8.7292545e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101110100010101010001010111000;
		b = 32'b01100110000110100010101111111110;
		correct = 32'b00000111111001100011001111001100;
		#400 //6.304418e-11 * 1.8201399e+23 = 3.4636997e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001100000100010100101011101110;
		b = 32'b10110001111001110111000101111010;
		correct = 32'b01011001101000001011010101101001;
		#400 //-38087610.0 * -6.7358856e-09 = 5654432400000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000000001101000010000110010000;
		b = 32'b01010011010010100010100111111001;
		correct = 32'b10101100011001000001100110001110;
		#400 //-2.8145485 * 868287600000.0 = -3.2414934e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110011111010101000110000001;
		b = 32'b00001111101111110001101011001000;
		correct = 32'b01101110001010011010101110010000;
		#400 //0.24738123 * 1.884437e-29 = 1.3127593e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111101001111001001011111111100;
		b = 32'b01100001000010111110101010011101;
		correct = 32'b01011011101011001000100000001110;
		#400 //1.5667751e+37 * 1.613127e+20 = 9.712658e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111110000101110000101010100110;
		b = 32'b01011110100101100100010001010010;
		correct = 32'b11011111000000001010100011110000;
		#400 //-5.019218e+37 * 5.413935e+18 = -9.270924e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010100111110100011110010000000;
		b = 32'b01001000100101111101001100101111;
		correct = 32'b01001011110100101111011111100011;
		#400 //8598055000000.0 * 310937.47 = 27652038.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101110111111101111100000001000;
		b = 32'b11010010011001001000000110010110;
		correct = 32'b11011100000011101101001011000110;
		#400 //3.9454522e+28 * -245356660000.0 = -1.6080478e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010101100110000001101000110010;
		b = 32'b01000001110100111000111101000101;
		correct = 32'b01010011001110000000110110010100;
		#400 //20904784000000.0 * 26.444956 = 790501800000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101011011100000010100000011101;
		b = 32'b11111101001100011000001000011100;
		correct = 32'b00101101101011010010110011100110;
		#400 //-2.9033163e+26 * -1.4746808e+37 = 1.9687762e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000101010010011010111100111;
		b = 32'b10000100001000011111001100111100;
		correct = 32'b01101100000001011011110100001000;
		#400 //-1.2311688e-09 * -1.9037147e-36 = 6.467192e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010000100111110001110011000000;
		b = 32'b10100101001110100011000111101100;
		correct = 32'b01101010110110101100001110010000;
		#400 //-21355692000.0 * -1.6149843e-16 = 1.3223467e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000100000011001110001101010100;
		b = 32'b00110101011010011111101011010101;
		correct = 32'b10001110000110100010010110101110;
		#400 //-1.6561305e-36 * 8.716427e-07 = -1.9000108e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011111111110110010100010010010;
		b = 32'b11100000000110101100111010100011;
		correct = 32'b10111111010011111010101010101001;
		#400 //3.6195751e+19 * -4.462013e+19 = -0.8111978
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000111000100010000110111100110;
		b = 32'b10010000001101011011011100100001;
		correct = 32'b00110110010011000101101000011110;
		#400 //-1.0912672e-34 * -3.5837033e-29 = 3.0450824e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010010011010100100110001001110;
		b = 32'b01000110001111000110101000010000;
		correct = 32'b10001011100111110010101111011011;
		#400 //-7.3931434e-28 * 12058.516 = -6.131056e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000101101111011011111100101110;
		b = 32'b11011010101010011000101000001110;
		correct = 32'b00101010100011110100000110100101;
		#400 //-6071.8975 * -2.3860532e+16 = 2.5447453e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100100010110010110010000111011;
		b = 32'b11011110100010001000011111111001;
		correct = 32'b01000101010010111100111011001110;
		#400 //-1.6040663e+22 * -4.919053e+18 = 3260.9253
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001000100010100101110011101011;
		b = 32'b00111110000001011001111010110110;
		correct = 32'b11001010000001001000101100100011;
		#400 //-283367.34 * 0.13048825 = -2171592.8
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100011001011000011000101010010;
		b = 32'b10101010110010100111010111001010;
		correct = 32'b01110111110110011011101001111010;
		#400 //-3.176394e+21 * -3.596414e-13 = 8.832114e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101001010010010010001101101110;
		b = 32'b00111111011000000001000000010010;
		correct = 32'b11101001011001011100111011011100;
		#400 //-1.5197588e+25 * 0.8752452 = -1.7363805e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101111111011110111110010111000;
		b = 32'b01000010001000000110111111101100;
		correct = 32'b00101101001111110001000101010010;
		#400 //4.3562465e-10 * 40.1093 = 1.0860939e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110001000011101100000001001000;
		b = 32'b10101001001111000101111101011110;
		correct = 32'b11000111010000100000000000000100;
		#400 //2.0773019e-09 * -4.1827104e-14 = -49664.016
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011101000001101001111101100010;
		b = 32'b01101101011101101110111011101010;
		correct = 32'b00101111000010111001000011001010;
		#400 //6.0628624e+17 * 4.776384e+27 = 1.2693416e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110101111111011001111001000111;
		b = 32'b11110011001100101011111011001001;
		correct = 32'b10000010001101011001110111100110;
		#400 //1.8896034e-06 * -1.4161658e+31 = -1.3343094e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101010110110001100111110000011;
		b = 32'b11000010110100100001000111001110;
		correct = 32'b00100111100001000001101110000011;
		#400 //-3.8513298e-13 * -105.034775 = 3.666719e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010011111010111110101000011011;
		b = 32'b01111101110001100101100111101110;
		correct = 32'b00010101100110000011110110000010;
		#400 //2026489900000.0 * 3.295676e+37 = 6.1489353e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100001000100000101011010010010;
		b = 32'b11000100010110010000101010011110;
		correct = 32'b11011100001010100011111100100000;
		#400 //1.6641057e+20 * -868.1659 = -1.9168061e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010011000001001110011001111010;
		b = 32'b01001011011100011010000011010101;
		correct = 32'b01000111000011001100111000010111;
		#400 //570802440000.0 * 15835349.0 = 36046.09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001111000000111010111010001101;
		b = 32'b01101000100101111110000000000001;
		correct = 32'b10100101110111011111011001100011;
		#400 //-2209254700.0 * 5.737676e+24 = -3.8504347e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101110010110101010010100100001;
		b = 32'b11101101001001001001100111100110;
		correct = 32'b00000000101010100000011011001010;
		#400 //-4.9714125e-11 * -3.1838496e+27 = 1.561447e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110011110100011010101101011100;
		b = 32'b11100011100001100111110101101000;
		correct = 32'b10001111110001111000110100111011;
		#400 //9.763491e-08 * -4.9618004e+21 = -1.9677315e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110011011100001110011011000101;
		b = 32'b01011010001101111111110111111010;
		correct = 32'b11011000101001111001011100111111;
		#400 //-1.9086179e+31 * 1.2947293e+16 = -1474144300000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101110001000001000010110011110;
		b = 32'b11011000110010000000000100011000;
		correct = 32'b11010100110011010111011010110101;
		#400 //1.2419784e+28 * -1759256200000000.0 = -7059679000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101110010110110110111110110000;
		b = 32'b11100111001011011000101000111101;
		correct = 32'b00000110101000011101101000101111;
		#400 //-4.9894033e-11 * -8.1951945e+23 = 6.088206e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101001010110100101111101100111;
		b = 32'b01000000111100101001010001011111;
		correct = 32'b00100111111001100111010000110001;
		#400 //4.8488472e-14 * 7.5806117 = 6.39638e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100011001101000110010111010111;
		b = 32'b11001101011111101011000000100110;
		correct = 32'b10010101001101010101001110111010;
		#400 //9.779385e-18 * -267059800.0 = -3.6618708e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000100000000100111010011110010;
		b = 32'b00100001111001110111110101001001;
		correct = 32'b10100001100100000100010100010110;
		#400 //-1.5335125e-36 * 1.5686332e-18 = -9.776106e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111000110100001010100111110100;
		b = 32'b11001010001011101011100110011100;
		correct = 32'b11101110000110001101110011100111;
		#400 //3.385765e+34 * -2862695.0 = -1.1827194e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111010011110100011011010101110;
		b = 32'b10001000111100111001010011000110;
		correct = 32'b11110001000000110111110000111101;
		#400 //0.0009544891 * -1.4660007e-33 = -6.510837e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000101001011010011100111101111;
		b = 32'b00101110101110111010100110111000;
		correct = 32'b10010101111011000100111001100111;
		#400 //-8.1450616e-36 * 8.5339236e-11 = -9.544334e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110001010000011011100111001111;
		b = 32'b00110110011001111101110101110000;
		correct = 32'b10111010010101011110010000010001;
		#400 //-2.8190816e-09 * 3.4550576e-06 = -0.000815929
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101010000001000010010001110101;
		b = 32'b11100010100100111010100111001111;
		correct = 32'b10000110111001010001011110000001;
		#400 //1.1736604e-13 * -1.3619537e+21 = -8.617476e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011011101101011010010110011101;
		b = 32'b01010000011110010011101111101010;
		correct = 32'b10001010101110101001001111111110;
		#400 //-3.0050963e-22 * 16725813000.0 = -1.7966817e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110111011000010101001100101101;
		b = 32'b01010011001000001011110111110000;
		correct = 32'b11100011101100110110110110001010;
		#400 //-4.570132e+33 * 690381400000.0 = -6.6197206e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101011010111101010001010011111;
		b = 32'b00010110111010001010110100011000;
		correct = 32'b01010011111101001111001111011100;
		#400 //7.9095926e-13 * 3.759086e-25 = 2104126600000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101111001100101010001000100101;
		b = 32'b10101110000011110100000110001010;
		correct = 32'b11000000100111111001110000100000;
		#400 //1.6246611e-10 * -3.2572646e-11 = -4.987808
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101010101010101011110000100000;
		b = 32'b01000010100100101010101110111001;
		correct = 32'b11100111100101010000000000110011;
		#400 //-1.0320289e+26 * 73.335396 = -1.4072726e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001010100000011101010000110101;
		b = 32'b01101010011010000011011101100011;
		correct = 32'b10011111100011110010000001000100;
		#400 //-4254234.5 * 7.0183087e+25 = -6.0616235e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011001001010010100111111111100;
		b = 32'b10011001011110110110100000100100;
		correct = 32'b11111111001011000110011111100001;
		#400 //2978576000000000.0 * -1.2997427e-23 = -2.2916659e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111100111100011010100010010010;
		b = 32'b01010011000000101001101100110110;
		correct = 32'b01101001011011001101011000001011;
		#400 //1.00381004e+37 * 560949760000.0 = 1.789483e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100011011001001110111011110110;
		b = 32'b11001101100010001110100011101101;
		correct = 32'b01010101010101100000100011101011;
		#400 //-4.2230766e+21 * -287120800.0 = 14708362000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101101000110010000000001000001;
		b = 32'b00010001110100001010000100001100;
		correct = 32'b11011010101110111011110110111000;
		#400 //-8.6970995e-12 * 3.2915866e-28 = -2.642221e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000011010011011100100111000101;
		b = 32'b11111101010111101100111000111011;
		correct = 32'b10000101011011000111001001111111;
		#400 //205.78816 * -1.8509964e+37 = -1.1117696e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100101111101110010001011100110;
		b = 32'b11000000010001101110101010111001;
		correct = 32'b01100101000111110000011101001010;
		#400 //-1.45883535e+23 * -3.1080763 = 4.693692e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000001110100100000011011001110;
		b = 32'b11001101101011110110100111101110;
		correct = 32'b10110011100110010100000111001111;
		#400 //26.253323 * -367869380.0 = -7.136588e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101100100000010011110011010011;
		b = 32'b01000110011101111011100111011110;
		correct = 32'b00100101100001011000110111011000;
		#400 //3.6731534e-12 * 15854.467 = 2.316794e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001111010001001100011111011000;
		b = 32'b00001111000101001101001100101010;
		correct = 32'b10111111101010010011111011010010;
		#400 //-9.7020346e-30 * 7.337632e-30 = -1.3222296
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011011110101000010110110110011;
		b = 32'b10100011110010110000011100011000;
		correct = 32'b01110111100001011100010011101001;
		#400 //-1.1944588e+17 * -2.2012308e-17 = 5.4263226e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011000001001100010000001010000;
		b = 32'b01101011010000101111011011100111;
		correct = 32'b00101100010110100010001000111000;
		#400 //730630850000000.0 * 2.3569757e+26 = 3.0998659e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110010101101101011001100101;
		b = 32'b11001001001000000000010110000000;
		correct = 32'b00101100101010111101100011001111;
		#400 //-3.201328e-06 * -655448.0 = 4.884183e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010100111011100011110111110;
		b = 32'b10110011100011000001101110001010;
		correct = 32'b01000110100100000010010100111101;
		#400 //-0.0012037677 * -6.524267e-08 = 18450.62
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101000010010101111110110101101;
		b = 32'b00111010111000110101000101001011;
		correct = 32'b01101100111001001001101010011000;
		#400 //3.83439e+24 * 0.0017342953 = 2.2109211e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011000101001100110111110001101;
		b = 32'b10111100010111000000010100111000;
		correct = 32'b01011011110000011010011100011010;
		#400 //-1463984300000000.0 * -0.013428979 = 1.090168e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101000110110000111101111111111;
		b = 32'b01101000110100011011101011001010;
		correct = 32'b00111111100001000001111101011010;
		#400 //8.178548e+24 * 7.923362e+24 = 1.0322068
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000100110001000111111101010010;
		b = 32'b10010011110110010011100001101001;
		correct = 32'b00110000011001111001001111001111;
		#400 //-4.6196304e-36 * -5.4834126e-27 = 8.424736e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111000100110100010111101010001;
		b = 32'b01001100100110110101011110010100;
		correct = 32'b11101011011111100001011111000101;
		#400 //-2.501792e+34 * 81444000.0 = -3.071794e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000010010101101000110000001111;
		b = 32'b01000011100100110010111000000000;
		correct = 32'b10111110001110101001011010100100;
		#400 //-53.636776 * 294.35938 = -0.18221527
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100001101011100111010010000000;
		b = 32'b01010000000001110011110100111001;
		correct = 32'b10010001001001010001110111100100;
		#400 //-1.1821536e-18 * 9075746000.0 = -1.3025416e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100100101111001100011010000001;
		b = 32'b11011000010111000111001000000100;
		correct = 32'b00001011110110110011100011011101;
		#400 //-8.186828e-17 * -969529000000000.0 = 8.444129e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010110100111001010111000010111;
		b = 32'b11010100110011111001100111000010;
		correct = 32'b10000001010000010011010100111100;
		#400 //2.5313025e-25 * -7133103000000.0 = -3.5486695e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111001011010001100000101010011;
		b = 32'b01000101001001000010000011000000;
		correct = 32'b11110011101101011000010101011111;
		#400 //-7.553337e+34 * 2626.0469 = -2.8763148e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111100011110010110101000100101;
		b = 32'b11011011110101010011000011100011;
		correct = 32'b00100000000101011011111110101100;
		#400 //-0.015223061 * -1.2001584e+17 = 1.268421e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110100011100001101101000101110;
		b = 32'b10111110101000111111111011010101;
		correct = 32'b11110101001110111111110011001100;
		#400 //7.632913e+31 * -0.3203036 = -2.3830245e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011001000100001111001100011110;
		b = 32'b10011110110000100111001100111010;
		correct = 32'b00111001101111101101010011000000;
		#400 //-7.493723e-24 * -2.0588206e-20 = 0.00036398135
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100111000001111011100100010111;
		b = 32'b10001101101111100011101011010001;
		correct = 32'b01011000101101101010010111100101;
		#400 //-1.883535e-15 * -1.1723814e-30 = 1606589000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010011110111001011010001100100;
		b = 32'b00111001101001011110001110010100;
		correct = 32'b11011001101010100100101110111001;
		#400 //-1895838500000.0 * 0.0003164081 = -5991750500000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010110100001101001101111110111;
		b = 32'b10111001011010010010001110110000;
		correct = 32'b00011100100100111100111011110100;
		#400 //-2.1747295e-25 * -0.00022233906 = 9.78114e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100001010001100010111101101100;
		b = 32'b11011000011100011101111011101110;
		correct = 32'b01001000010100011100001100110010;
		#400 //-2.2849203e+20 * -1063759100000000.0 = 214796.78
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011001010110111010101000101101;
		b = 32'b00010010000101001101100110101000;
		correct = 32'b01000110101111001110010100101010;
		#400 //1.1356401e-23 * 4.696885e-28 = 24178.582
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100001100000011100001110100100;
		b = 32'b10000110110011100101001011011000;
		correct = 32'b11011010001000010000000111101001;
		#400 //8.793166e-19 * -7.7610316e-35 = -1.1329893e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111001111011000000111101000100;
		b = 32'b00110000011101010100011111001000;
		correct = 32'b11001000111101100110000001010010;
		#400 //-0.00045024802 * 8.923249e-10 = -504578.56
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100001111100010010011110010101;
		b = 32'b10010010100000111110010101011100;
		correct = 32'b01001110111010100000100000001010;
		#400 //-1.6341272e-18 * -8.323804e-28 = 1963197700.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001010010101001101010110010010;
		b = 32'b01111000110101000111011001101000;
		correct = 32'b00010001000000000011100101010101;
		#400 //3487076.5 * 3.4474016e+34 = 1.0115086e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100000010110100111010100111110;
		b = 32'b10100010011110111001111001010110;
		correct = 32'b11111101010111100100001100010101;
		#400 //6.2966225e+19 * -3.4100666e-18 = -1.8464808e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111000111011101101101100011001;
		b = 32'b01000001001010000010000000000101;
		correct = 32'b01110111001101011101100110011011;
		#400 //3.8756578e+34 * 10.507817 = 3.6883566e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000110010111011011100110000010;
		b = 32'b00000010010001111111100101000001;
		correct = 32'b01000011100011011110110000100111;
		#400 //4.170177e-35 * 1.4691743e-37 = 283.84494
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001001111010001000010110000101;
		b = 32'b10101111000010111101111001101111;
		correct = 32'b00011010010101001100101001011010;
		#400 //-5.597753e-33 * -1.2721e-10 = 4.400403e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100101000010011001100101011000;
		b = 32'b11111000100100101001110000111010;
		correct = 32'b00101011111100000100001111100100;
		#400 //-4.0612056e+22 * -2.3788875e+34 = 1.7071869e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110101000111001100000010011011;
		b = 32'b11001111100100100000001011011110;
		correct = 32'b10100101000010010110101010001011;
		#400 //5.8394807e-07 * -4899323000.0 = -1.1918954e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011001001001011010101110011011;
		b = 32'b11101101101101001111011011000100;
		correct = 32'b00101010111010100101110101101111;
		#400 //-2914503300000000.0 * -7.000703e+27 = 4.1631583e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000011000001100000100111010011;
		b = 32'b11101000110111000100110000111000;
		correct = 32'b10011001100110111100001011011010;
		#400 //134.03838 * -8.322613e+24 = -1.6105324e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000110100000010110011000100011;
		b = 32'b00000000110111111110011001000111;
		correct = 32'b11000101000100111111001101101111;
		#400 //-4.8674483e-35 * 2.0561924e-38 = -2367.2146
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001100010100001101110100001101;
		b = 32'b11110100110000001001111111001100;
		correct = 32'b00010111000010101100101010000101;
		#400 //-54752308.0 * -1.220901e+32 = 4.484582e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110000001000001000110001000111;
		b = 32'b10001010100011001111110001010001;
		correct = 32'b01100101000100011100001010110011;
		#400 //-5.8407007e-10 * -1.357642e-32 = 4.302092e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011011110011110011100101111110;
		b = 32'b01100100101110101010111110101111;
		correct = 32'b00110110100011100001010011111010;
		#400 //1.1665707e+17 * 2.755003e+22 = 4.2343718e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100110111011100000001010111100;
		b = 32'b00001000100011010001111100001000;
		correct = 32'b01011101110101111110000101111111;
		#400 //1.6515309e-15 * 8.493424e-34 = 1.9444818e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100100010001001000101000010000;
		b = 32'b01001100100101111000110010110010;
		correct = 32'b01010111001001011111111110101001;
		#400 //1.4502041e+22 * 79455630.0 = 182517470000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101110011100101110000000111011;
		b = 32'b10010010101101000000100110010000;
		correct = 32'b01011011001011001010110100001001;
		#400 //-5.5223586e-11 * -1.1361954e-27 = 4.860395e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010011110001011001101111101;
		b = 32'b01000001111100011100110010011100;
		correct = 32'b10111000000000111010011101010011;
		#400 //-0.0009487195 * 30.224907 = -3.1388667e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110011001011000011011111101111;
		b = 32'b00111111001101111001010010100101;
		correct = 32'b11110011011100000010011111011010;
		#400 //-1.3644555e+31 * 0.7171119 = -1.9027092e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101110011100111011010010111100;
		b = 32'b01011110111101101010010010011101;
		correct = 32'b10001110111111001111001110011001;
		#400 //-5.5412328e-11 * 8.8862513e+18 = -6.2357372e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000001010100111010101100100001;
		b = 32'b11011000010001001111011010111111;
		correct = 32'b00101000100010011000111001011000;
		#400 //-13.2292795 * -866256200000000.0 = 1.5271787e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101011101010101100110111111011;
		b = 32'b00110011110011111000100010011000;
		correct = 32'b10110111010100101011000110001011;
		#400 //-1.2136398e-12 * 9.664035e-08 = -1.2558313e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110101010000101110010011001;
		b = 32'b10011001010010100001011010000101;
		correct = 32'b01011100110101010100011011000011;
		#400 //-5.01757e-06 * -1.0447703e-23 = 4.802558e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001001010010010011000011000011;
		b = 32'b01011001100011110000011010111110;
		correct = 32'b00101111001101000000110110101101;
		#400 //824076.2 * 5032292000000000.0 = 1.6375763e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101000101000100111010000011111;
		b = 32'b00011011111110100110010111000101;
		correct = 32'b01001100001001100001011010100000;
		#400 //1.8035972e-14 * 4.1424798e-22 = 43539070.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110111011011000111001000100110;
		b = 32'b11010010011110010001000111000101;
		correct = 32'b11100100011100110000011001110101;
		#400 //4.7956924e+33 * -267436240000.0 = -1.7932096e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010010000000100000011010000101;
		b = 32'b01000011000000011100111110000000;
		correct = 32'b10001110100000000011011001000001;
		#400 //-4.1028803e-28 * 129.81055 = -3.160668e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001010000001001110000101110011;
		b = 32'b10101101100111100100100100011101;
		correct = 32'b00011011110101101110100101101110;
		#400 //-6.397971e-33 * -1.799499e-11 = 3.555418e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111111110010001000010010101000;
		b = 32'b11111100100101000001100001100000;
		correct = 32'b10000010101011010100111101000100;
		#400 //1.5665483 * -6.1516346e+36 = -2.5465562e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010100110010011111100001100111;
		b = 32'b10100000000011101010001101100010;
		correct = 32'b00110100001101010011111001000000;
		#400 //-2.0393791e-26 * -1.2081927e-19 = 1.6879585e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111101110001010001100111101001;
		b = 32'b11100001110100011101111011111101;
		correct = 32'b00011011011100000110110001100100;
		#400 //-0.096240826 * -4.839297e+20 = 1.9887358e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001001101011101110011100101000;
		b = 32'b10011100100010100111100100000100;
		correct = 32'b11101100101000011010110011001110;
		#400 //1432805.0 * -9.163356e-22 = -1.5636248e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110010000110000110010110101001;
		b = 32'b10111111110110011101001011110001;
		correct = 32'b01110001101100110001101100111010;
		#400 //-3.0185357e+30 * -1.7017499 = 1.7737834e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111100001010011000101010011;
		b = 32'b11100100001000001000110000000011;
		correct = 32'b10100010110101000110000111011110;
		#400 //68194.65 * -1.1846272e+22 = -5.7566336e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000010110011001010000110001010;
		b = 32'b10110000001011011011101101100110;
		correct = 32'b00010010000101101100001111101110;
		#400 //-3.0067825e-37 * -6.320334e-10 = 4.7573156e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011111001101110100001110101011;
		b = 32'b10110111100110001001111000011111;
		correct = 32'b11100111000110011011010000001010;
		#400 //1.3205587e+19 * -1.8193443e-05 = -7.258432e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001101110100110010100001110101;
		b = 32'b00111110000100111110110110100011;
		correct = 32'b11001111001101101011011000110011;
		#400 //-442830500.0 * 0.1444612 = -3065394000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100100101010011000110111101110;
		b = 32'b10101111110011101101011111111001;
		correct = 32'b11110100010100011101100101010111;
		#400 //2.5021815e+22 * -3.762464e-10 = -6.6503798e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101111000101000000110110000110;
		b = 32'b11010011111011110111101111110010;
		correct = 32'b11011010100111100100001101011111;
		#400 //4.582013e+28 * -2057153300000.0 = -2.227356e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010101100101010101001110000010;
		b = 32'b00101110010101110000110111111000;
		correct = 32'b01100110101100011100000111011011;
		#400 //20523237000000.0 * 4.8897747e-11 = 4.1971743e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010100101001110000110010111110;
		b = 32'b10100011000001000011101101110111;
		correct = 32'b11110001001000011011001111111111;
		#400 //5739786500000.0 * -7.1683265e-18 = -8.00715e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101001101100100101111000001010;
		b = 32'b11100110100111001100100100010000;
		correct = 32'b00000010100100011001111010011011;
		#400 //-7.921101e-14 * -3.7019906e+23 = 2.139687e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001001010001001000001101000011;
		b = 32'b00000001100001101110100001001001;
		correct = 32'b11000111001110100111001101111101;
		#400 //-2.365436e-33 * 4.955714e-38 = -47731.49
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011110111110011001011010101;
		b = 32'b11010010000111100100001011100110;
		correct = 32'b00111001001101001000010101000001;
		#400 //-29255082.0 * -169931800000.0 = 0.00017215779
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011001011001111100101001000110;
		b = 32'b11101011110001101110100111010100;
		correct = 32'b10101101000101010010011111110011;
		#400 //4077695000000000.0 * -4.8094307e+26 = -8.47854e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100101011100101001011101011001;
		b = 32'b11101111110010100000010001011111;
		correct = 32'b10110101000110011011010101001010;
		#400 //7.1600285e+22 * -1.2504251e+29 = -5.726075e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000011011111000000111110011101;
		b = 32'b11111011100000011110101001111001;
		correct = 32'b10000111011110000101100000000001;
		#400 //252.06099 * -1.349124e+36 = -1.8683308e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100100011001001100110010110100;
		b = 32'b11100010110011011001101010010111;
		correct = 32'b11000001000011100111000011001111;
		#400 //1.6882432e+22 * -1.896361e+21 = -8.902541
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011110000011001010000001110100;
		b = 32'b01011111010010111101000001111001;
		correct = 32'b00111110001100001010001000110001;
		#400 //2.5333067e+18 * 1.4686371e+19 = 0.17249371
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010110101100110111010111010001;
		b = 32'b11101110110001101001001000100010;
		correct = 32'b00100111011001110101110011000100;
		#400 //-98659300000000.0 * -3.0727348e+28 = 3.2107978e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000110100110001110010010100101;
		b = 32'b10011010110100001001001110101100;
		correct = 32'b11101011001110111010011111011111;
		#400 //19570.322 * -8.626536e-23 = -2.2686188e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101101011100111111000101110100;
		b = 32'b11110001110100100110000011011101;
		correct = 32'b00111011000101000110101111111000;
		#400 //-4.7185473e+27 * -2.0834865e+30 = 0.0022647362
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111110101110111010000111011000;
		b = 32'b11110011100101111000110010110010;
		correct = 32'b11001010100111100111100111000101;
		#400 //1.2470299e+38 * -2.4013991e+31 = -5192930.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011011011011101110000110111000;
		b = 32'b10101101000000000111001111011000;
		correct = 32'b10101101111011100000101001001001;
		#400 //1.9759832e-22 * -7.30168e-12 = -2.7062035e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101010000000011100101000101111;
		b = 32'b11011000001100111101100000110010;
		correct = 32'b11010001001110001011111111011111;
		#400 //3.9226554e+25 * -790964500000000.0 = -49593315000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110101110110110011011000010011;
		b = 32'b11101010000101111000011010010000;
		correct = 32'b01001011001110010010110101000101;
		#400 //-5.557665e+32 * -4.5795813e+25 = 12135749.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110100100001110010011110011010;
		b = 32'b10010000110110101010001111000010;
		correct = 32'b01100011000111100011111111011010;
		#400 //-2.5174523e-07 * -8.623815e-29 = 2.9191866e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011010110110010001010001010000;
		b = 32'b11100110100101101110010001011011;
		correct = 32'b00110011101110000010010101011110;
		#400 //-3.0551202e+16 * -3.562837e+23 = 8.574965e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000111011001000000100011010001;
		b = 32'b00010111010011111100110100110110;
		correct = 32'b00101111100011000111011001111110;
		#400 //1.7155404e-34 * 6.714432e-25 = 2.5550045e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000111011110110011011000100100;
		b = 32'b00001110000101111000110101101011;
		correct = 32'b00111000110101000010101111011001;
		#400 //1.8899052e-34 * 1.8680277e-30 = 0.00010117115
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111010100010010101111001011001;
		b = 32'b01100101100111111110011000111001;
		correct = 32'b00010100010110111110110110010111;
		#400 //0.0010480388 * 9.438789e+22 = 1.1103531e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000010000101011101101000010101;
		b = 32'b01101100111100011010000110000011;
		correct = 32'b00010100100111101100001101011101;
		#400 //37.46297 * 2.3369107e+27 = 1.603098e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000000110111110111010111011101;
		b = 32'b10101000000011010010101000101011;
		correct = 32'b01011000010010101001111011111000;
		#400 //-6.9831376 * -7.836216e-15 = 891136460000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011101001000000011101110011100;
		b = 32'b11110111101100111100001111110011;
		correct = 32'b10100100111001000010111100100000;
		#400 //7.216246e+17 * -7.292152e+33 = -9.895907e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001111101001011011001101011001;
		b = 32'b10101001111111110100111011100101;
		correct = 32'b10100101001001100010011001001011;
		#400 //1.6339338e-29 * -1.1337961e-13 = -1.4411179e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110100110111000110010011000101;
		b = 32'b10101101001010011100011111110000;
		correct = 32'b11000111001001100010100001010001;
		#400 //4.1051513e-07 * -9.650933e-12 = -42536.316
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100001001110101001010101100010;
		b = 32'b10000110111001011001100111010001;
		correct = 32'b01011001110100000000100101100000;
		#400 //-6.321696e-19 * -8.636624e-35 = 7319638000000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111100100001001000000110110100;
		b = 32'b00111111100111001111001111110110;
		correct = 32'b11111100010110000010000001100101;
		#400 //-5.504111e+36 * 1.2261951 = -4.4887726e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111111100101100110101101000101;
		b = 32'b01101010100101111101110001000001;
		correct = 32'b10010100011111011001000111111011;
		#400 //-1.1751486 * 9.179396e+25 = -1.2802025e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100100100011101100101011001001;
		b = 32'b00111100110010111111010100101011;
		correct = 32'b01100111001100110011101000110000;
		#400 //2.10724e+22 * 0.024897179 = 8.46377e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011101100000011011100110001000;
		b = 32'b10100110100001101010101010111111;
		correct = 32'b10110110011101101001101011011000;
		#400 //3.433785e-21 * -9.344399e-16 = -3.6746987e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110010111011000101101101001001;
		b = 32'b10100000000110001111000101101000;
		correct = 32'b11010010010001011100111101010111;
		#400 //2.7515528e-08 * -1.2954775e-19 = -212396790000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001110011101011011100111100011;
		b = 32'b10011000011110100111110010010011;
		correct = 32'b11110101011110110010001001111101;
		#400 //1030650050.0 * -3.2374637e-24 = -3.1835108e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110000011010011011101101100;
		b = 32'b11100000000100010010101010111010;
		correct = 32'b10011101011110010000100010010100;
		#400 //0.13790673 * -4.184151e+19 = -3.295931e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110001111010010010101111010001;
		b = 32'b10111001100100100100100011000101;
		correct = 32'b01110111110011000000011011011100;
		#400 //-2.3092153e+30 * -0.00027901508 = 8.27631e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001101010010100111010100000001;
		b = 32'b00110000111110100101110111111100;
		correct = 32'b11011011110011110000001100010100;
		#400 //-212291600.0 * 1.8216606e-09 = -1.1653741e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011110111100010101010110001101;
		b = 32'b00110001001100101110110100110101;
		correct = 32'b11101101001011001010010100011101;
		#400 //-8.6949803e+18 * 2.6037246e-09 = -3.3394395e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101011110011101010111110001100;
		b = 32'b11001101001100101100100001110101;
		correct = 32'b01011110000100111111101000011011;
		#400 //-4.9973543e+26 * -187467600.0 = 2.6657162e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010100001110000110001110101011;
		b = 32'b00010010100010111011101001010001;
		correct = 32'b01000001001010001110100110110111;
		#400 //9.309282e-27 * 8.818064e-28 = 10.557059
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110100110100001010000001110001;
		b = 32'b11010001000110010000110010110001;
		correct = 32'b10100011001011100111101100011001;
		#400 //3.8859756e-07 * -41083933000.0 = -9.458626e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110011000111111010101010101000;
		b = 32'b00110010111010011011001100010111;
		correct = 32'b10111111101011101110011100001111;
		#400 //-3.7175283e-08 * 2.720621e-08 = -1.3664263
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100111001010101001101010101011;
		b = 32'b10111000110000101110100110011110;
		correct = 32'b00101101111000000001001010111000;
		#400 //-2.3676085e-15 * -9.2941555e-05 = 2.5474164e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110001110010101100110111111000;
		b = 32'b00000011111011100110010000011011;
		correct = 32'b11101101010110011100100011101111;
		#400 //-5.9023897e-09 * 1.4011366e-36 = -4.2125726e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011100000001100010001010101011;
		b = 32'b10010001010100001100001110101100;
		correct = 32'b11001010001001000111110000111101;
		#400 //4.438169e-22 * -1.6468603e-28 = -2694927.2
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110100000010110100110011111110;
		b = 32'b11100111010111010111000100000010;
		correct = 32'b10001100001000010000101001010000;
		#400 //1.2973393e-07 * -1.0457276e+24 = -1.2406092e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111000001111011010111010111101;
		b = 32'b01001100111000111010010010100110;
		correct = 32'b01101010110101010100111110001111;
		#400 //1.5388878e+34 * 119350580.0 = 1.2893845e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101001111100011001101010001111;
		b = 32'b11111111001011101111111011101110;
		correct = 32'b10101010001100001011100001011001;
		#400 //3.6510126e+25 * -2.3260934e+38 = -1.5695899e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000101100110000010011101000110;
		b = 32'b10100111001000111000111111010011;
		correct = 32'b00011101111011100010010011100001;
		#400 //-1.4308438e-35 * -2.2698761e-15 = 6.3036207e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011101010001101110001110001101;
		b = 32'b10001111010000111010101111111100;
		correct = 32'b11001101100000100001101010111110;
		#400 //2.6322723e-21 * -9.647365e-30 = -272848830.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011101110101110011100000101001;
		b = 32'b11000111111001001001001111011001;
		correct = 32'b10010101011100010000101000001101;
		#400 //5.6968094e-21 * -117031.695 = -4.867749e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011000011000001000011110001001;
		b = 32'b00100111001101010110000011001101;
		correct = 32'b01110000100111100111001111000101;
		#400 //987490900000000.0 * 2.5171272e-15 = 3.923087e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001100100000101100100100111101;
		b = 32'b10001101100110000100011010110000;
		correct = 32'b10111110010110111101111100110100;
		#400 //2.0150787e-31 * -9.384741e-31 = -0.21471864
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000000101000100101001011111010;
		b = 32'b10001111111110011010111100000101;
		correct = 32'b01110000001001100110111000110101;
		#400 //-5.072629 * -2.462071e-29 = 2.0603098e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100011000000010100011110010110;
		b = 32'b00111001001101100011111110101011;
		correct = 32'b00101001001101011001100010000010;
		#400 //7.008263e-18 * 0.0001738059 = 4.0322353e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000000011011101001000100001101;
		b = 32'b10001111001001100111100110001001;
		correct = 32'b01110000101101110110111000101101;
		#400 //-3.7276032 * -8.207839e-30 = 4.541516e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110010001000001010010011000110;
		b = 32'b10100011010100101010111100110100;
		correct = 32'b11001110010000110011001000110100;
		#400 //9.350691e-09 * -1.14212235e-17 = -818711800.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001000111111100110100000001101;
		b = 32'b01101110001010001100100110010101;
		correct = 32'b00011010010000001110110111100001;
		#400 //521024.4 * 1.3059295e+28 = 3.9896826e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100000100110000011111000011110;
		b = 32'b00001001001101010101111001100101;
		correct = 32'b11010110110101101110001110001100;
		#400 //-2.5790907e-19 * 2.1831467e-33 = -118136400000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101100011111011101100011100001;
		b = 32'b10100111100101110001010001111011;
		correct = 32'b11000100010101110001000101011010;
		#400 //3.6073854e-12 * -4.1933124e-15 = -860.2711
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111100110010010111000101011101;
		b = 32'b01000001100010010011111011001101;
		correct = 32'b10111010101110111101111101111001;
		#400 //-0.024590189 * 17.155664 = -0.0014333568
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010100011110111111110100101010;
		b = 32'b10110111101001111110011001111101;
		correct = 32'b11011100010000000001101100000011;
		#400 //4329136700000.0 * -2.001528e-05 = -2.1629158e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110111010011101001101001101010;
		b = 32'b11000110101001010010010111111100;
		correct = 32'b11110000001000000010000101000111;
		#400 //4.1904103e+33 * -21138.992 = -1.9823133e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111010011010001110010100011110;
		b = 32'b11101101101111101111001110001011;
		correct = 32'b10001100000111000001110110110010;
		#400 //0.0008884239 * -7.387072e+27 = -1.2026739e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101000101010101000011100100100;
		b = 32'b01011001101101111110001000100011;
		correct = 32'b01001110011011010110100000011110;
		#400 //6.4423617e+24 * 6469820000000000.0 = 995755900.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111001110001110100010100001001;
		b = 32'b01100100101000110010111100001001;
		correct = 32'b01010100100111000100111000110110;
		#400 //1.2933341e+35 * 2.4081668e+22 = 5370616500000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101111100110011110110010011001;
		b = 32'b01111101110101001110110011111011;
		correct = 32'b00110001001110010001000000001011;
		#400 //9.527447e+28 * 3.537835e+37 = 2.6930163e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010000100101101101100100010111;
		b = 32'b10001111000000001001010011111100;
		correct = 32'b01000001000101100010101001001110;
		#400 //-5.949905e-29 * -6.3395806e-30 = 9.385328
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001011100100111111100111010101;
		b = 32'b11100110101101000000011110110011;
		correct = 32'b10100100010100100110101101100010;
		#400 //19395498.0 * -4.25084e+23 = -4.5627448e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100101010011111001111100100001;
		b = 32'b01011100000110100010000111101001;
		correct = 32'b11001000101011000110101110011000;
		#400 //-6.127908e+22 * 1.7353772e+17 = -353116.75
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100011011110110011000101100101;
		b = 32'b01011110101011111100111001101111;
		correct = 32'b10000100001101101110001100010001;
		#400 //-1.3617197e-17 * 6.3340924e+18 = -2.1498261e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100111011001101011111001000001;
		b = 32'b10100011011000000100110000000100;
		correct = 32'b01000011100000111010110110111111;
		#400 //-3.2022049e-15 * -1.2159161e-17 = 263.3574
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110010110001011000101100000111;
		b = 32'b11011010111101101001101010001110;
		correct = 32'b10010111010011010001000111101100;
		#400 //2.299704e-08 * -3.470639e+16 = -6.6261693e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000001111100011001101000110000;
		b = 32'b00011010001101110111000000111010;
		correct = 32'b01100111001010001001010111110010;
		#400 //30.200287 * 3.793417e-23 = 7.961236e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111101101101111111101000011000;
		b = 32'b11110110000100001010010011000100;
		correct = 32'b01000111001000101100111010110000;
		#400 //-3.056841e+37 * -7.334303e+32 = 41678.688
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010010110001001010001110010000;
		b = 32'b10111100101100111011101010001000;
		correct = 32'b00010101100011000000101100010010;
		#400 //-1.240966e-27 * -0.021939531 = 5.6563016e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101110000111001111101010111110;
		b = 32'b11010100010010101010100110101010;
		correct = 32'b10011001010001100100101100101110;
		#400 //3.5692997e-11 * -3481719500000.0 = -1.02515425e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001000111010010011110001100110;
		b = 32'b01001010101110111001000001001001;
		correct = 32'b00111101100111110010101100011100;
		#400 //477667.2 * 6146084.5 = 0.07771894
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100010100010101101011111011000;
		b = 32'b11000100000000101000101011110010;
		correct = 32'b10011110000010000010001110000010;
		#400 //3.763351e-18 * -522.171 = -7.207123e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110101001101001011000101101111;
		b = 32'b10000100101000010010100010011101;
		correct = 32'b11110000000011111000001111100101;
		#400 //6.7313425e-07 * -3.7888216e-36 = -1.7766323e+29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110010101110001011100111010110;
		b = 32'b11110101011010110000110001001101;
		correct = 32'b10111100110010010011000100110100;
		#400 //7.3177477e+30 * -2.979588e+32 = -0.024559595
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001010110011001010111111000001;
		b = 32'b10010100111011011111010111010000;
		correct = 32'b00110101010111000011010000110000;
		#400 //-1.9710597e-32 * -2.402784e-26 = 8.203233e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100010100011111110101101100010;
		b = 32'b10010101001000110010001101011100;
		correct = 32'b11001100111000011101011101110110;
		#400 //3.900945e-18 * -3.294548e-26 = -118406060.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011011010111001001100110111000;
		b = 32'b01110100011100011110010010100100;
		correct = 32'b10100110011010010111011100110000;
		#400 //-6.209351e+16 * 7.665899e+31 = -8.0999643e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011011110101011100101100001001;
		b = 32'b01010100110101000110011111001011;
		correct = 32'b00000110100000001101011000010100;
		#400 //3.5369102e-22 * 7298195400000.0 = 4.846281e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001111110001000001111111101100;
		b = 32'b10010011000100010000111001111110;
		correct = 32'b00111100001011010001000000101110;
		#400 //-1.9339388e-29 * -1.8308718e-27 = 0.01056294
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111111101001000001101100101010;
		b = 32'b11110100100001110111001101111010;
		correct = 32'b10001010100110110001010000101000;
		#400 //1.282079 * -8.585232e+31 = -1.4933539e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001110110100111010011000101001;
		b = 32'b01001001100000001100011111001011;
		correct = 32'b11000100110100100101110111001110;
		#400 //-1775441000.0 * 1054969.4 = -1682.9314
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000010011111110001100110001111;
		b = 32'b11011011100011010001101011100010;
		correct = 32'b10100110011001110110100001011100;
		#400 //63.77496 * -7.943506e+16 = -8.028566e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111100100000011000100011011101;
		b = 32'b10101010011111011110110110100110;
		correct = 32'b01010001100000101001011101101000;
		#400 //-0.015812332 * -2.2553365e-13 = 70110740000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111011011100000010010110001001;
		b = 32'b01000100111110101110101101001011;
		correct = 32'b01110101111101010000001001100110;
		#400 //1.24691255e+36 * 2007.3529 = 6.2117255e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101011000101100000001100000001;
		b = 32'b01111100101111101111010100011101;
		correct = 32'b00101101110010010001101110001101;
		#400 //1.8135306e+26 * 7.932063e+36 = 2.286329e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101110100101001001001001011111;
		b = 32'b11001100010110101110100110010010;
		correct = 32'b10100001101011011011111000010000;
		#400 //6.7562615e-11 * -57386570.0 = -1.1773245e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000000001101101111000000101000;
		b = 32'b11010010000000001110000010111111;
		correct = 32'b00101101101101011011000100100011;
		#400 //-2.858408 * -138381600000.0 = 2.0655982e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100000000010100001010110111110;
		b = 32'b10101101110011011001001000111011;
		correct = 32'b10110001101010111111010101101000;
		#400 //1.1696249e-19 * -2.3370741e-11 = -5.0046545e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101001001001001001000100011001;
		b = 32'b01111100010011111001001010110011;
		correct = 32'b00101100010010101111010111011010;
		#400 //1.2434315e+25 * 4.3111235e+36 = 2.8842402e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000100010111010010110101110010;
		b = 32'b10001101110110000011111010010011;
		correct = 32'b10110110000000101110101110000110;
		#400 //2.5999293e-36 * -1.3327092e-30 = -1.9508602e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001101110001110001011110010011;
		b = 32'b11101011011001111000100011101000;
		correct = 32'b00100001110111000010000100010101;
		#400 //-417526370.0 * -2.7990839e+26 = 1.4916537e-18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110100011011110111000000101110;
		b = 32'b01100000111111100010110111111101;
		correct = 32'b10010010111100010010011100101010;
		#400 //-2.229942e-07 * 1.4652459e+20 = -1.5218893e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011101001110111000000110010110;
		b = 32'b10100001111111110111101000111101;
		correct = 32'b01111010101110111110001111000010;
		#400 //-8.444528e+17 * -1.7311828e-18 = 4.877895e+35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011110011001111110100011111011;
		b = 32'b11011001110000010001100001100000;
		correct = 32'b00000100000110011011101011010101;
		#400 //-1.22772174e-20 * -6793934000000000.0 = 1.8070853e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111010101110110000101001101110;
		b = 32'b01010001100101010110001011100110;
		correct = 32'b10101000101000000100001110000110;
		#400 //-0.0014270076 * 80201170000.0 = -1.7792852e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000100010100000000100111011111;
		b = 32'b00100100101110110011110101101011;
		correct = 32'b11011111000011100011011111100000;
		#400 //-832.15424 * 8.120237e-17 = -1.0247906e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000101010110011010011110001110;
		b = 32'b00001111011001111110011101100010;
		correct = 32'b10110101011100000100010100100100;
		#400 //-1.0234066e-35 * 1.1433742e-29 = -8.950758e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110011011000010000001001001101;
		b = 32'b11101101110001011001001000000010;
		correct = 32'b00000101000100011100011011010101;
		#400 //-5.2388987e-08 * -7.6431324e+27 = 6.854387e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100101110111101101001011110011;
		b = 32'b01000010000100000010101100101001;
		correct = 32'b01100011010001011101010110001100;
		#400 //1.3153209e+23 * 36.04215 = 3.6493963e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010110011011111111010111011100;
		b = 32'b11001100011011001110010000001110;
		correct = 32'b01001001100000011010100010011001;
		#400 //-65959810000000.0 * -62099510.0 = 1062163.1
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111111001111110101010011111100;
		b = 32'b11010100011110111110111110110000;
		correct = 32'b01101010010000100110101100001100;
		#400 //-2.5432381e+38 * -4328232300000.0 = 5.875928e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000001101110110100101001111000;
		b = 32'b10001001101010001001010100110000;
		correct = 32'b00110111100011100011010001011101;
		#400 //-6.879981e-38 * -4.0584824e-33 = 1.6952103e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000011100101011110111000011111;
		b = 32'b10100110000111110010101100110110;
		correct = 32'b11011100111100010010010000011000;
		#400 //299.86032 * -5.522277e-16 = -5.4300124e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001101000110001100010110000110;
		b = 32'b11001011110011000000110000101100;
		correct = 32'b11000000101111111010101100101110;
		#400 //160192600.0 * -26744920.0 = -5.989646
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010000110100001001001011111011;
		b = 32'b10010001011000110011101110101110;
		correct = 32'b01111110111010101111101010010111;
		#400 //-27994348000.0 * -1.7925533e-28 = 1.5617024e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111111011110000010011001011001;
		b = 32'b11000000001111000010000000110111;
		correct = 32'b10111110101010001101011100001101;
		#400 //0.96933514 * -2.9394662 = -0.3297657
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010011110100011100011010111001;
		b = 32'b11000111001110111011111101111010;
		correct = 32'b10001100000011110000010010100100;
		#400 //5.2954973e-27 * -48063.477 = -1.1017716e-31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001010111111001100001111100001;
		b = 32'b01000101110111000111100001000110;
		correct = 32'b00000100100100101011111111111110;
		#400 //2.4340399e-32 * 7055.034 = 3.4500752e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000010101011100010111111001101;
		b = 32'b00110000110000010000001110101011;
		correct = 32'b00010001011001110000011101001000;
		#400 //2.5594438e-37 * 1.4043641e-09 = 1.8224931e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110000110101001001000101011000;
		b = 32'b10110011010100011111011100010000;
		correct = 32'b10111101000000011001011000101111;
		#400 //1.5466339e-09 * -4.8886307e-08 = -0.031637367
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001011010110000101100111010110;
		b = 32'b00011010011001100000100110011000;
		correct = 32'b10110000011100001100010011001101;
		#400 //-4.1667672e-32 * 4.7570635e-23 = -8.759116e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000000010100010011100110101101;
		b = 32'b01100000110000001110111000111111;
		correct = 32'b00011111000010101100111110001010;
		#400 //3.2691453 * 1.1121695e+20 = 2.939431e-20
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000101110110000001101011000001;
		b = 32'b01110100011010011000000011011001;
		correct = 32'b00010000111011001110110011001000;
		#400 //6915.344 * 7.4000153e+31 = 9.3450406e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010010100110000011001100100100;
		b = 32'b11010001000110110110001000011110;
		correct = 32'b00000000111110101100000101001011;
		#400 //-9.605156e-28 * -41710380000.0 = 2.3028214e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101010111101001101000011111011;
		b = 32'b10011010111111100110001111001000;
		correct = 32'b11001111011101100101110110110000;
		#400 //4.3488116e-13 * -1.0521314e-22 = -4133335000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110110000010001101111010111000;
		b = 32'b11100010011110100000001111001100;
		correct = 32'b10010011000011000010010110000101;
		#400 //2.0395219e-06 * -1.1529899e+21 = -1.7688983e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001001100101001111001001010100;
		b = 32'b01111010011111111001000001010000;
		correct = 32'b00001110100101010011001101101100;
		#400 //1220170.5 * 3.3174068e+35 = 3.6780853e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100110011110100111000110000111;
		b = 32'b00110111101110000111100010010001;
		correct = 32'b10101110001011011100011011011001;
		#400 //-8.689003e-16 * 2.1990652e-05 = -3.9512258e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011011000000010000101001110001;
		b = 32'b01111111010010110000011000111100;
		correct = 32'b00011011001000101011011000110011;
		#400 //3.6321752e+16 * 2.6986565e+38 = 1.3459198e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110011111001101110010000101001;
		b = 32'b00001010000000000101101101100000;
		correct = 32'b01101001011001100011111111001011;
		#400 //1.0751712e-07 * 6.1801615e-33 = 1.7397137e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111010100101101111100011101011;
		b = 32'b00101100111101100100011110100111;
		correct = 32'b01001101000111001110111001001110;
		#400 //0.0011518275 * 6.9996955e-12 = 164553950.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011110000011111011100101000111;
		b = 32'b11011011011110000011100000010001;
		correct = 32'b00000010000101000011101010100101;
		#400 //-7.6086714e-21 * -6.986744e+16 = 1.0890153e-37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110111000011100100111111000010;
		b = 32'b10011111011101011001101111111011;
		correct = 32'b11010111000101000101010100001000;
		#400 //8.48243e-06 * -5.2009792e-20 = -163092930000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001001101100010101111001101011;
		b = 32'b00111001100111000001111001010100;
		correct = 32'b00001111100100010110110001000111;
		#400 //4.269999e-33 * 0.00029777235 = 1.4339811e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111110010001110011100111011111;
		b = 32'b01010001111111000001100011010100;
		correct = 32'b11101011110010100100111101111110;
		#400 //-6.6204214e+37 * 135343540000.0 = -4.891568e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000010100000111000101111001100;
		b = 32'b10010101010111000010000111011001;
		correct = 32'b00101100100110001111101011011000;
		#400 //-1.932896e-37 * -4.4455347e-26 = 4.347949e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010001000001011001010100110001;
		b = 32'b10100010011010110101110110101111;
		correct = 32'b00101110000100010100101100110000;
		#400 //-1.0537823e-28 * -3.1898034e-18 = 3.3035963e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111101110110001111100001110000;
		b = 32'b10010101111000011101111100000101;
		correct = 32'b11100111011101011110100101111011;
		#400 //0.10594261 * -9.122864e-26 = -1.16128674e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111101000001011111010001110000;
		b = 32'b10101010010010000111000010110001;
		correct = 32'b11010010001010110001010111101100;
		#400 //0.032703817 * -1.7802666e-13 = -183701800000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100001101110101110111110011100;
		b = 32'b00110110110110011110001001000001;
		correct = 32'b01101010010110111010001101100010;
		#400 //4.31045e+20 * 6.4934434e-06 = 6.6381577e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010011110100111001010101010111;
		b = 32'b00100100001100111101111010101010;
		correct = 32'b11101111000101101001000101110110;
		#400 //-1817487200000.0 * 3.900304e-17 = -4.6598603e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000010011000001100011010011100;
		b = 32'b00000101011110011101011110000100;
		correct = 32'b11111100011001100101000011101110;
		#400 //-56.193954 * 1.1747508e-35 = -4.783479e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000011000000000000000101111011;
		b = 32'b00100111000110001001110011111101;
		correct = 32'b11011011010101101011100011101111;
		#400 //-128.00578 * 2.117934e-15 = -6.043898e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110110100100101000101110111011;
		b = 32'b01101111111010111011111100100001;
		correct = 32'b11000110000111110010001011000110;
		#400 //-1.4861512e+33 * 1.4592008e+29 = -10184.693
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001110111111001111101010100111;
		b = 32'b10001000000001111011101001100010;
		correct = 32'b01000110011011101001001100110110;
		#400 //-6.2364166e-30 * -4.0844177e-34 = 15268.803
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101100100101111000011000000100;
		b = 32'b01011100100101100101110001100011;
		correct = 32'b00001111100000001111110101011110;
		#400 //4.306557e-12 * 3.385826e+17 = 1.2719368e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000001110111010100101100111110;
		b = 32'b10000100101111000111010111110101;
		correct = 32'b11111100100101100100110011000001;
		#400 //27.66174 * -4.4306914e-36 = -6.24321e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011111010011101111000111100100;
		b = 32'b01010111010011011001101000110110;
		correct = 32'b01000111100000001101010111110110;
		#400 //1.491195e+19 * 226062210000000.0 = 65963.92
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101101001101101111011110001110;
		b = 32'b10011010000100010000100001100001;
		correct = 32'b01010010101000010111101010110001;
		#400 //-1.040047e-11 * -2.9992066e-23 = 346774080000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011110001010111110100011101111;
		b = 32'b10011011101010011000100010111001;
		correct = 32'b01000010000000011100101100110101;
		#400 //-9.100834e-21 * -2.804706e-22 = 32.448444
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010101000011111001111001011010;
		b = 32'b11100101110010111101000010100110;
		correct = 32'b00101110101101000110010000001010;
		#400 //-9869392000000.0 * -1.2031116e+23 = 8.203223e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001011111000101100111010100110;
		b = 32'b10010011111010101111100110000011;
		correct = 32'b00110111011101110001101000001100;
		#400 //-8.7362963e-32 * -5.9315942e-27 = 1.4728412e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100100101000100000010100101110;
		b = 32'b11011000011101100101010011101101;
		correct = 32'b11001011101010000110000100011101;
		#400 //2.3909966e+22 * -1083378460000000.0 = -22069818.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100010101110110000100111001110;
		b = 32'b11100110111110001010110001010101;
		correct = 32'b00111011010000001000110010010100;
		#400 //-1.7251238e+21 * -5.8716293e+23 = 0.0029380666
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011010111000000101100110010100;
		b = 32'b11011001110001011111011010001010;
		correct = 32'b11000000100100010000111110110110;
		#400 //3.1574443e+16 * -6965205400000000.0 = -4.533168
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000001111000010001111000010111;
		b = 32'b11101111010001110001110000110011;
		correct = 32'b10010010000100001011100000011000;
		#400 //28.139692 * -6.162161e+28 = -4.56653e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000010010100011100111000001000;
		b = 32'b11011110001011100010111000010001;
		correct = 32'b00100011100110100010111000000010;
		#400 //-52.451202 * -3.137747e+18 = 1.6716199e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101100100001000001101010010100;
		b = 32'b11001111100111000010100110000111;
		correct = 32'b11011100010110001000111110000001;
		#400 //1.2776298e+27 * -5239934500.0 = -2.4382552e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011001111000100111110100000011;
		b = 32'b00110000001110110110101000100110;
		correct = 32'b11101001000110101010111110111011;
		#400 //-7968849600000000.0 * 6.818105e-10 = -1.1687777e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010000100111111100000100011111;
		b = 32'b10100011110111011010111101110111;
		correct = 32'b11101100001110000111101110010010;
		#400 //21441870000.0 * -2.403518e-17 = -8.921036e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100110011011110100111101101001;
		b = 32'b01010111101000000000011000011001;
		correct = 32'b10001110001111110110101101101111;
		#400 //-8.3027403e-16 * 351896100000000.0 = -2.3594295e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100111010110011101010111000010;
		b = 32'b11100101000001110010111010110101;
		correct = 32'b10000001110011100100001011010111;
		#400 //3.0230678e-15 * -3.9898817e+22 = -7.576836e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101111101010110110001011101110;
		b = 32'b00001110110000011110110101011100;
		correct = 32'b11100000011000100011111010001110;
		#400 //-3.1175013e-10 * 4.7806742e-30 = -6.5210495e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100011001000010111011010011000;
		b = 32'b01111000010000110011001100001011;
		correct = 32'b00101010010100111100000101111001;
		#400 //2.9784714e+21 * 1.5836456e+34 = 1.8807689e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101100111100110001111000011100;
		b = 32'b10010111011011011101001001111010;
		correct = 32'b01010101000000101101100110100000;
		#400 //-6.909818e-12 * -7.684449e-25 = 8991950000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100101001101010010001000100001;
		b = 32'b11001011010100100011001101000110;
		correct = 32'b00011001010111001001100110001001;
		#400 //-1.5710811e-16 * -13775686.0 = 1.14047396e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001010111001101001100010010100;
		b = 32'b01110011000100110110010111110101;
		correct = 32'b10010111010010000011111110100001;
		#400 //-7556170.0 * 1.1678094e+31 = -6.4703796e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010111101111100010111011110001;
		b = 32'b00100001010111100100001010011101;
		correct = 32'b10110101110110110000110111000101;
		#400 //-1.2290312e-24 * 7.530469e-19 = -1.6320779e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110111101010101111111100000001;
		b = 32'b00001100010010010110010101110000;
		correct = 32'b01101010110110010101101110001100;
		#400 //2.0384325e-05 * 1.5515002e-31 = 1.3138461e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110111011011111001001010000100;
		b = 32'b10101100110100010011000011110100;
		correct = 32'b11001010000100101001011011110000;
		#400 //1.4279623e-05 * -5.945572e-12 = -2401724.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001111111010100100000000001011;
		b = 32'b11011111100010001110010000011000;
		correct = 32'b10101111110110110000100100100111;
		#400 //7860131300.0 * -1.972807e+19 = -3.984237e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010100110011001101100110110000;
		b = 32'b01100110010111100101111001010000;
		correct = 32'b00101101111010111101010100011100;
		#400 //7038604000000.0 * 2.6252628e+23 = 2.6811046e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001010011101000110011101000011;
		b = 32'b00000110011000110010111110111010;
		correct = 32'b01000011100010011011001101000100;
		#400 //1.1767594e-32 * 4.272902e-35 = 275.4005
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001111001000011001100000001010;
		b = 32'b01111100101111110101101011001000;
		correct = 32'b00010001110110000010111101101010;
		#400 //2711095800.0 * 7.94856e+36 = 3.4108012e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110011001111101100110011000001;
		b = 32'b01110000110101111011001101001100;
		correct = 32'b01000001111000100111001001111110;
		#400 //1.5116719e+31 * 5.3404827e+29 = 28.305904
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010010111010101110100111010101;
		b = 32'b10111101101001100110001000100010;
		correct = 32'b01010100101101001011100010000001;
		#400 //-504472700000.0 * -0.08124186 = 6209516600000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100101011001010101110101110000;
		b = 32'b01100000010111100100100011111110;
		correct = 32'b11000100100001000001001110101100;
		#400 //-6.7696596e+22 * 6.4069325e+19 = -1056.6147
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010111010000010110011101010010;
		b = 32'b10110010111100101001011111111110;
		correct = 32'b10100011110011000001011101101110;
		#400 //6.249207e-25 * -2.8241626e-08 = -2.2127647e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000110110101011110100100111111;
		b = 32'b00011000010000110110011000010110;
		correct = 32'b11101110000011000010000001111100;
		#400 //-27380.623 * 2.52547e-24 = -1.0841793e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011110110010000100100100101011;
		b = 32'b00101110101101101110000111000100;
		correct = 32'b11101111100011000010111001011100;
		#400 //-7.216057e+18 * 8.316506e-11 = -8.676789e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111110010100001000100010010110;
		b = 32'b01001111100000010101111111111011;
		correct = 32'b10101110010011100101000100111111;
		#400 //-0.20364603 * 4341102000.0 = -4.6911138e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011010010100100101100101011010;
		b = 32'b11010000001100010010110111111000;
		correct = 32'b10001001100101111111011001110000;
		#400 //4.349916e-23 * -11890319000.0 = -3.6583676e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111000110110111111111110010011;
		b = 32'b00001010101011001100111010001010;
		correct = 32'b01101101101000101111010010010000;
		#400 //0.00010490338 * 1.6640689e-32 = 6.3040287e+27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001111100101010100000001011101;
		b = 32'b11100010000011011100101000110010;
		correct = 32'b10101101000001101011110001100101;
		#400 //5008046600.0 * -6.5389016e+20 = -7.65885e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011110111011010110100000101100;
		b = 32'b10100101011110101111100001101011;
		correct = 32'b01111000111100100010101000101011;
		#400 //-8.553486e+18 * -2.1768211e-16 = 3.9293472e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110100101010110010010111110011;
		b = 32'b01001111111010110000111011100010;
		correct = 32'b00100100001110100110010101101111;
		#400 //3.1878844e-07 * 7887242000.0 = 4.041824e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111101011111001010001111100100;
		b = 32'b01111011000100001011110000111100;
		correct = 32'b01000001110111110110110110011110;
		#400 //2.0988526e+37 * 7.515086e+35 = 27.928524
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111000111000100010010111101011;
		b = 32'b11101011010110000111011010000011;
		correct = 32'b01001101000001011011101000100011;
		#400 //-3.669463e+34 * -2.6168763e+26 = 140223020.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010111110111011010100111001000;
		b = 32'b01010000111101001010111000110110;
		correct = 32'b01000110011001111110101011111001;
		#400 //487442550000000.0 * 32840462000.0 = 14842.743
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011010110000100100011110110101;
		b = 32'b10010011101110101111000000101011;
		correct = 32'b11000110100001010000011011110100;
		#400 //8.035237e-23 * -4.7189825e-27 = -17027.477
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110111101011101100010000101111;
		b = 32'b11010000001000101100000110100001;
		correct = 32'b00100111000010010111000111111101;
		#400 //-2.0833771e-05 * -10922395000.0 = 1.9074362e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011110100100010000011011001100;
		b = 32'b11100110101001101101000101001100;
		correct = 32'b00110111010111101000111100101101;
		#400 //-5.225132e+18 * -3.9388684e+23 = 1.3265567e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111011010011001001100010011001;
		b = 32'b11001011010100001000001101001110;
		correct = 32'b00101111011110110011000011101111;
		#400 //-0.0031218885 * -13665102.0 = 2.2845702e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011010110011001101101110100;
		b = 32'b11111001000001100111000010001111;
		correct = 32'b00010001110011110010111100001111;
		#400 //-14261108.0 * -4.362817e+34 = 3.2687844e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110011000111000011001011101100;
		b = 32'b11010111100001101100111000110111;
		correct = 32'b11011011000101000101000000111001;
		#400 //1.2375353e+31 * -296440500000000.0 = -4.1746502e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101100010001100000001010011100;
		b = 32'b10001011001011101001001011010101;
		correct = 32'b01100000100100010010111100100001;
		#400 //-2.813894e-12 * -3.3621645e-32 = 8.369293e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100011100101110111110100101100;
		b = 32'b10000101101010101101011101011001;
		correct = 32'b01011101011000110000000001010100;
		#400 //-1.6424465e-17 * -1.606583e-35 = 1.0223229e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010001011100011011011000001001;
		b = 32'b11100001101101101110100001010011;
		correct = 32'b00101111001010010010011010110010;
		#400 //-64883823000.0 * -4.2175602e+20 = 1.5384208e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101011100100111111100111010001;
		b = 32'b10010111010100101001010010111010;
		correct = 32'b11010011101100111110010001010110;
		#400 //1.0514316e-12 * -6.804238e-25 = -1545260000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111100011010111000100101111111;
		b = 32'b11000010111001000011010011101011;
		correct = 32'b10111001000001000001110010010000;
		#400 //0.014376043 * -114.103355 = -0.00012599141
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011110101011111001111011110001;
		b = 32'b10110000101100001000001110100001;
		correct = 32'b00101101011111101011010001010101;
		#400 //-1.8594582e-20 * -1.2843097e-09 = 1.447827e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101001110010100100000111111100;
		b = 32'b01110011110110000010011010100001;
		correct = 32'b00110101011011111000101110101001;
		#400 //3.0564327e+25 * 3.4250476e+31 = 8.923767e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011101100010111100011111001101;
		b = 32'b00110101011100001101100010100001;
		correct = 32'b01100111100101001001001101001000;
		#400 //1.2590306e+18 * 8.9722204e-07 = 1.4032542e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110010111000100010101001011111;
		b = 32'b01011011111011111000000100100101;
		correct = 32'b10010110011100011011111000001010;
		#400 //-2.632913e-08 * 1.3482903e+17 = -1.9527791e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000011000101101101011110101001;
		b = 32'b10110001101010001101100011101001;
		correct = 32'b01010000111001001011001110100000;
		#400 //-150.84242 * -4.9141033e-09 = 30695817000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101000010111110110011000111110;
		b = 32'b00111100011011010101001101011000;
		correct = 32'b00101011011100001111101001011111;
		#400 //1.2401157e-14 * 0.014485203 = 8.561259e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100001100010110010000101101011;
		b = 32'b00010101111111100110001011101011;
		correct = 32'b01001011000011000000001101011000;
		#400 //9.427852e-19 * 1.0274585e-25 = 9175896.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11101011011110100101001001110101;
		b = 32'b11010100010010101001110100110000;
		correct = 32'b01010110100111100010001110100110;
		#400 //-3.0262085e+26 * -3480882200000.0 = 86937970000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111000001011000000110000101111;
		b = 32'b01001111110110000010010101000001;
		correct = 32'b01100111110010111100010101011111;
		#400 //1.3958159e+34 * 7252640300.0 = 1.9245625e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010100101000101101000011100111;
		b = 32'b00000100001110010011001001111011;
		correct = 32'b01001111111000010000111111110010;
		#400 //1.6440217e-26 * 2.1769825e-36 = 7551837000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000100001111000001110010111011;
		b = 32'b00011010000100110011001111110101;
		correct = 32'b11101001101000111001001010010100;
		#400 //-752.4489 * 3.0440858e-23 = -2.4718388e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001100111100110010111111110011;
		b = 32'b10010000010111001000000001001011;
		correct = 32'b01111100000011010010101101010010;
		#400 //-127500184.0 * -4.3486183e-29 = 2.93197e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010100000001110100110001101101;
		b = 32'b01100111100110001001110000010100;
		correct = 32'b10101011111000101111010111111100;
		#400 //-2324411200000.0 * 1.4413577e+24 = -1.612654e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001101011100111101110110001111;
		b = 32'b11010000111001000100010100110010;
		correct = 32'b00111100000010001011111010101100;
		#400 //-255711470.0 * -30637920000.0 = 0.008346241
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011010101000101001111010000101;
		b = 32'b10011011000111111011010100111010;
		correct = 32'b10111111000000100101010101010011;
		#400 //6.725773e-23 * -1.3210729e-22 = -0.50911444
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010110100101010010000011101000;
		b = 32'b11001101111000010110111100111101;
		correct = 32'b00001000001010010101100100011100;
		#400 //-2.4093015e-25 * -472770460.0 = 5.0961335e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011010011001111111001010100011;
		b = 32'b00101110100000011100100010110001;
		correct = 32'b00101011011001001100001001110010;
		#400 //4.796568e-23 * 5.901891e-11 = 8.127172e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101011101000100110111000101100;
		b = 32'b10011000001100111100101010110000;
		correct = 32'b11010010111001110100011110010111;
		#400 //1.1541371e-12 * -2.3237539e-24 = -496669260000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011011101011010101101110000101;
		b = 32'b00110010110011100110000001000011;
		correct = 32'b01101000010101110000101011000011;
		#400 //9.7591596e+16 * 2.4025331e-08 = 4.0620292e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010110111000101101000111001101;
		b = 32'b11000010111000001110001100100111;
		correct = 32'b00010011100000010001100110001010;
		#400 //-3.6644672e-25 * -112.44366 = 3.258936e-27
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100101010000110111101011101100;
		b = 32'b00101011000101001101101100100100;
		correct = 32'b00111001101010000001011101111010;
		#400 //1.6955201e-16 * 5.288428e-13 = 0.00032060948
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100000011010001111110110011110;
		b = 32'b01101011000010010010010111110100;
		correct = 32'b00110100110110010111001100001101;
		#400 //6.7154995e+19 * 1.6580207e+26 = 4.050311e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110110000100011110110000111101;
		b = 32'b00111110101111010110101111100101;
		correct = 32'b01110110110001010011011001011000;
		#400 //7.399165e+32 * 0.3699638 = 1.9999701e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110001011110001001101111000100;
		b = 32'b01100010011001001100110110000100;
		correct = 32'b10001110100010110001010001111000;
		#400 //-3.6177292e-09 * 1.05516665e+21 = -3.4285856e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110111001000111101000101101100;
		b = 32'b01001000000011111111110100000011;
		correct = 32'b01101110100100011010000010111011;
		#400 //3.322625e+33 * 147444.05 = 2.2534819e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011000100001101101110001110111;
		b = 32'b01010000101101100101110101100101;
		correct = 32'b11000111001111010101000010111100;
		#400 //-1186251600000000.0 * 24476592000.0 = -48464.734
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010010000111101111010000010000;
		b = 32'b00101000101010001110010010111001;
		correct = 32'b00101000111100001110111011101111;
		#400 //5.015684e-28 * 1.875094e-14 = 2.6748974e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000000000110010111011011100111;
		b = 32'b11111001110111011100110100111111;
		correct = 32'b10000101101100010010000001001111;
		#400 //2.3978822 * -1.4395756e+35 = -1.6656868e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100000100100001111101010111100;
		b = 32'b01111001101011101110101110101111;
		correct = 32'b10100110010101000010111000110000;
		#400 //-8.357495e+19 * 1.1352999e+35 = -7.361487e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100101111111110111011110011;
		b = 32'b01011110110111010010100100100101;
		correct = 32'b00100101010111100010101100100100;
		#400 //1535.4672 * 7.9681547e+18 = 1.9270047e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111111110000110110011010110000;
		b = 32'b11111100111001001010001001100100;
		correct = 32'b11111111110000110110011010110000;
		#400 //nan * -9.497099e+36 = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000001101010011110110010010011;
		b = 32'b00111001111001001111110010010001;
		correct = 32'b00000111001111011111100001010000;
		#400 //6.242026e-38 * 0.00043675725 = 1.4291752e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000000000001000101000001100001;
		b = 32'b00011000011011100010011111010110;
		correct = 32'b00100101000101000110010000010010;
		#400 //3.96177e-40 * 3.0780891e-24 = 1.2870859e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101011010000111001011000001110;
		b = 32'b10010000010011000100101100110001;
		correct = 32'b01011010011101010001011010101100;
		#400 //-6.948616e-13 * -4.0289832e-29 = 1.7246574e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111110111111000110000001101011;
		b = 32'b11110100101111000010110010000101;
		correct = 32'b01001001101010111010110000001111;
		#400 //-1.6773304e+38 * -1.1926938e+32 = 1406337.9
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101100011100010111100010111110;
		b = 32'b00101011110010011111101011101110;
		correct = 32'b11000000000110010000011011011001;
		#400 //-3.4315185e-12 * 1.4351556e-12 = -2.391043
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000000101111010100111010000010;
		b = 32'b10010101100110101100010101111100;
		correct = 32'b01101010100111001000111111000010;
		#400 //-5.9158335 * -6.251168e-26 = 9.463565e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001010011001000000101111010001;
		b = 32'b01000011001111101111101000101000;
		correct = 32'b01000110100110001101100001010011;
		#400 //3736308.2 * 190.97717 = 19564.162
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011111001011101111111110100101;
		b = 32'b01111010111110011001111100100011;
		correct = 32'b00100011101100110111100001011111;
		#400 //1.2609979e+19 * 6.480548e+35 = 1.9458198e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111110000010110110010001101000;
		b = 32'b10000100000101100011010101011111;
		correct = 32'b01111001011011011001000011011100;
		#400 //-0.1361252 * -1.7656922e-36 = 7.709453e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001000111001111001101000011101;
		b = 32'b11101000001010110001100111101101;
		correct = 32'b10100000001011010100001010100011;
		#400 //474320.9 * -3.2320117e+24 = -1.4675718e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110101000011011001011110011000;
		b = 32'b01100001011011100011110011010110;
		correct = 32'b01010011000110000010011000011110;
		#400 //1.794894e+32 * 2.746693e+20 = 653474500000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001100101011110111101010111000;
		b = 32'b11010011101001001111110101101110;
		correct = 32'b00111000100010000010001101000011;
		#400 //-92001730.0 * -1417253000000.0 = 6.491553e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010000100101111110100100000010;
		b = 32'b10101000000101000010110110001100;
		correct = 32'b01101000000000110011100101011010;
		#400 //-20389040000.0 * -8.225527e-15 = 2.4787518e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000001111110110110111101111100;
		b = 32'b10011010100001111010000100100001;
		correct = 32'b00100110111011010100101010110001;
		#400 //-9.236281e-38 * -5.609501e-23 = 1.6465424e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100101111011100010010001101001;
		b = 32'b01100010001010011000111111110011;
		correct = 32'b01000011001100111100010100011011;
		#400 //1.4057436e+23 * 7.819681e+20 = 179.76994
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100010110010100101011001101010;
		b = 32'b00011100111110001101111100001010;
		correct = 32'b11000101010100000010001000100101;
		#400 //-5.4843704e-18 * 1.6468918e-21 = -3330.134
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111011001101101110111101111000;
		b = 32'b11000110000110110011000111010111;
		correct = 32'b01110100100101101110000100110111;
		#400 //-9.49855e+35 * -9932.46 = 9.56314e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111100001110010100111001011010;
		b = 32'b11100101101010111011000100100111;
		correct = 32'b11010110000010100010011001001010;
		#400 //3.8486563e+36 * -1.0134907e+23 = -37974264000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111101100000000101101111001110;
		b = 32'b00001000100010101110000011100100;
		correct = 32'b11110100011011001001101110111011;
		#400 //-0.0626751 * 8.358444e-34 = -7.498417e+31
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11111101101100110010011001000100;
		b = 32'b11110110100110110110111000111001;
		correct = 32'b01000110100100111000100001110001;
		#400 //-2.9766312e+37 * -1.5762531e+33 = 18884.22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101011111000000010001000000001;
		b = 32'b01011000110101000011010011100010;
		correct = 32'b01010010100001110011000110011001;
		#400 //5.4191993e+26 * 1866588800000000.0 = 290326350000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110111001101101011101100001;
		b = 32'b10001010010111110010011010010111;
		correct = 32'b01101100000001000110100101001110;
		#400 //-6.8796076e-06 * -1.07443174e-32 = 6.40302e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010100110011010111000000101110;
		b = 32'b10001101111101110000111001011100;
		correct = 32'b11000110010101001110000000011110;
		#400 //2.0743957e-26 * -1.5226007e-30 = -13624.029
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000111010100000000110011011001;
		b = 32'b10101101111010011110000000110100;
		correct = 32'b00011000111000111011101100111001;
		#400 //-1.5651956e-34 * -2.65886e-11 = 5.886717e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011011111111100110011110001000;
		b = 32'b10010001100011001001010111011011;
		correct = 32'b01001001111001111010000100111100;
		#400 //-4.208768e-22 * -2.218046e-28 = 1897511.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100000111101001111100100111000;
		b = 32'b01110010100011101011010000001011;
		correct = 32'b00101101110110111011101110100000;
		#400 //1.4121761e+20 * 5.65306e+30 = 2.498074e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011111100010011001100011001010;
		b = 32'b01010101011001111110010001000110;
		correct = 32'b00001001100101111110011011100011;
		#400 //5.8274525e-20 * 15935476000000.0 = 3.6569053e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111100110001000011011010000101;
		b = 32'b00000000011111010100000001000000;
		correct = 32'b01111011110010001000010011111100;
		#400 //0.023951778 * 1.1502486e-38 = 2.0823132e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100001011101001000111111001011;
		b = 32'b11100001110011001001111010000101;
		correct = 32'b10111111000110001111110001110001;
		#400 //2.8196043e+20 * -4.718198e+20 = -0.59760195
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110110000001101011100101011100;
		b = 32'b11001011100100111101111100100101;
		correct = 32'b00101001111010010011110100001100;
		#400 //-2.007545e-06 * -19381834.0 = 1.03578685e-13
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11110111000100101101110011001110;
		b = 32'b11100000001010010011111110011001;
		correct = 32'b01010110010111100010001111000111;
		#400 //-2.9787258e+33 * -4.878254e+19 = 61061310000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011000000101100101100100111000;
		b = 32'b10111100110110001001010110010011;
		correct = 32'b01011010101100011011010111001011;
		#400 //-661239740000000.0 * -0.02643851 = 2.5010477e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110110101010011100001001000110;
		b = 32'b00010110101111100110010001100111;
		correct = 32'b01011111011001000100000110110000;
		#400 //5.059209e-06 * 3.0759518e-25 = 1.6447621e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000101101000101011010001101000;
		b = 32'b00111010010010000000011000100101;
		correct = 32'b10001010110100000011110010101111;
		#400 //-1.5300678e-35 * 0.000763031 = -2.0052498e-32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000100110100011100100010111110;
		b = 32'b01001110100001100010101010111011;
		correct = 32'b10110101110010000010010000111011;
		#400 //-1678.2732 * 1125473700.0 = -1.4911706e-06
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010010001010101111010010101101;
		b = 32'b11111001011011110011110100011101;
		correct = 32'b10011000001101101110111011011110;
		#400 //183562350000.0 * -7.7637405e+34 = -2.3643546e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101110111110000111010110001010;
		b = 32'b11110000100011000111010001011101;
		correct = 32'b10111101111000100110110101110000;
		#400 //3.844719e+28 * -3.477486e+29 = -0.1105603
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00000001111011111000100100101111;
		b = 32'b10010111110111111001000001110110;
		correct = 32'b10101001100010010010010011110111;
		#400 //8.7991583e-38 * -1.4447504e-24 = -6.0904346e-14
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011000010000011101001010111101;
		b = 32'b01110100011011101001011011011111;
		correct = 32'b00100011010011111111011110010101;
		#400 //852443400000000.0 * 7.561198e+31 = 1.127392e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100011001001111000101111101101;
		b = 32'b11111110110001110001111001110000;
		correct = 32'b00100011110101110110100010011011;
		#400 //-3.090689e+21 * -1.3233721e+38 = 2.3354649e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001101010011000110100111110110;
		b = 32'b11000010000110010111111000010010;
		correct = 32'b01001010101010100111011011011010;
		#400 //-214343520.0 * -38.373116 = 5585773.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010111100010001110101100011011;
		b = 32'b10110001001010110100001011110001;
		correct = 32'b10100101110011001010101000001101;
		#400 //8.848143e-25 * -2.4921827e-09 = -3.550359e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100000110011010101101001100000;
		b = 32'b00111000000111000001001101111010;
		correct = 32'b01101000001010000110100110100100;
		#400 //1.1837796e+20 * 3.7211437e-05 = 3.1812252e+24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111011100000101110000100011110;
		b = 32'b01111001101101000011111101000000;
		correct = 32'b01000001001110011110001001101000;
		#400 //1.359129e+36 * 1.1698704e+35 = 11.617775
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110110111100011110111100101001;
		b = 32'b01110001001010000000010100011100;
		correct = 32'b00000101001110000100111100010111;
		#400 //7.2102016e-06 * 8.319945e+29 = 8.666165e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110110111101001011001111011011;
		b = 32'b00000000011011101010000100001110;
		correct = 32'b01110110000011011001000000010001;
		#400 //7.2927046e-06 * 1.015968e-38 = 7.178085e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010110100101111100101001000001;
		b = 32'b11101000110000010011010110001011;
		correct = 32'b00101101010010010001111011000010;
		#400 //-83447465000000.0 * -7.2992354e+24 = 1.1432357e-11
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011100001000100101001010010001;
		b = 32'b10111100110001001110111011010111;
		correct = 32'b11011110110100110000001000111001;
		#400 //1.8275892e+17 * -0.024039669 = -7.602389e+18
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101101010111111100101010101001;
		b = 32'b00101010011011010010101011100110;
		correct = 32'b11000010011100011000111111011100;
		#400 //-1.2721082e-11 * 2.1064712e-13 = -60.390488
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010110111001101011111001000110;
		b = 32'b10110001011001000111001100010111;
		correct = 32'b10100101000000010100100100000000;
		#400 //3.7278584e-25 * -3.3243788e-09 = -1.12137e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001010000001111110101000100010;
		b = 32'b00010101001111001000100101000111;
		correct = 32'b00110100001110001000110001111101;
		#400 //6.544049e-33 * 3.807459e-26 = 1.7187445e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010000101111011111001111010101;
		b = 32'b11001010100000010010101001100001;
		correct = 32'b00000101101111000011110100001000;
		#400 //-7.492304e-29 * -4232496.5 = 1.7701854e-35
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001111101011000101000111000111;
		b = 32'b10011110111010111010110110001001;
		correct = 32'b10110000001110110010110110100011;
		#400 //1.6992009e-29 * -2.4953365e-20 = -6.809506e-10
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110010010010110110100010010110;
		b = 32'b10001100110111100001000001000000;
		correct = 32'b11100100111010100111111010000001;
		#400 //1.1839935e-08 * -3.4214296e-31 = -3.460523e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110000110011000101010100110100;
		b = 32'b01100111111100100111110001010111;
		correct = 32'b00001000010101111011100010000101;
		#400 //1.486717e-09 * 2.2902127e+24 = 6.491611e-34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10001000111010010010001110011101;
		b = 32'b11000100011011001010001010010000;
		correct = 32'b00000011111111000011011111010000;
		#400 //-1.403155e-33 * -946.54004 = 1.4824043e-36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011111011111100111101011010111;
		b = 32'b11001000110000111110010110000011;
		correct = 32'b01010110001001100100011101011001;
		#400 //-1.8337205e+19 * -401196.1 = 45706340000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011010011011111010000000111011;
		b = 32'b00101000101011110100111011010001;
		correct = 32'b00110001001011101111011000100000;
		#400 //4.9553475e-23 * 1.9463084e-14 = 2.5460238e-09
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011011100111000010100100101011;
		b = 32'b11000010111001110001111100101110;
		correct = 32'b00011000001011001111100001011011;
		#400 //-2.583464e-22 * -115.5609 = 2.2355866e-24
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111110010101010011100000001000;
		b = 32'b01000000000000011100000000010011;
		correct = 32'b10111101110100100101011110110110;
		#400 //-0.20822155 * 2.0273483 = -0.10270636
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011011000010000101101001010110;
		b = 32'b10001000000000100011011001000100;
		correct = 32'b11010010100001100000100101011101;
		#400 //1.1278845e-22 * -3.918424e-34 = -287841350000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111110011001010110000110011110;
		b = 32'b00111001100011010011001100011101;
		correct = 32'b01000100010011111111000000110000;
		#400 //0.22400519 * 0.00026931698 = 831.7529
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000110011110111111110010101001;
		b = 32'b11101010000101011100110101111111;
		correct = 32'b10011011110101110100111111100010;
		#400 //16127.165 * -4.5275094e+25 = -3.562039e-22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100100001100011110011111011010;
		b = 32'b11000000001011011000011100011011;
		correct = 32'b01100011100000110011101010110011;
		#400 //-1.3127121e+22 * -2.7113712 = 4.8415064e+21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011101010001001010111010101111;
		b = 32'b01110111000100111100010010010001;
		correct = 32'b00100101101010100101111011110100;
		#400 //8.857786e+17 * 2.9970878e+33 = 2.9554642e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100111001100111010010001111001;
		b = 32'b11010100011110100111001011001101;
		correct = 32'b01010010001101111001111111100000;
		#400 //-8.483376e+23 * -4302671400000.0 = 197165320000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011001001000010100101001111111;
		b = 32'b11010010100000000100101111011101;
		correct = 32'b01000110001000001110101100011111;
		#400 //-2837461300000000.0 * -275514300000.0 = 10298.78
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110011101100101000100110001111;
		b = 32'b11001110111100101010111100101001;
		correct = 32'b10100100001111000101010101011110;
		#400 //8.313793e-08 * -2035782800.0 = -4.083831e-17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001110010101001110111101001011;
		b = 32'b11111111111011101110011110100101;
		correct = 32'b11111111111011101110011110100101;
		#400 //-893113000.0 * nan = nan
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000111001111010001000110001010;
		b = 32'b10011010111010000000011001010010;
		correct = 32'b11101011110100001001101011101001;
		#400 //48401.54 * -9.596316e-23 = -5.0437623e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10011111000010111011010001100101;
		b = 32'b11000100011110010110011010000000;
		correct = 32'b00011010000011110110011011001010;
		#400 //-2.9583614e-20 * -997.60156 = 2.965474e-23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001011001010100101110010001101;
		b = 32'b10010011101010001010010100101011;
		correct = 32'b01110111000000010100110101111101;
		#400 //-11164813.0 * -4.257203e-27 = 2.62257e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000101000001110100111101011111;
		b = 32'b11100011101110010000110010000110;
		correct = 32'b10100000101110110011000010111010;
		#400 //2164.9607 * -6.8271e+21 = -3.1711277e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101101100000011111110111101111;
		b = 32'b11011100010111110111110011001000;
		correct = 32'b00010000100101001110011100100111;
		#400 //-1.4778371e-11 * -2.5162447e+17 = 5.8731854e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100000000100111000100010100010;
		b = 32'b11010111111110000011001011010010;
		correct = 32'b11000111100110000010101111001011;
		#400 //4.25237e+19 * -545794300000000.0 = -77911.586
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000001101010001100000010110100;
		b = 32'b01001001101000110111000111010100;
		correct = 32'b10110111100001000010100000110000;
		#400 //-21.094093 * 1338938.5 = -1.575434e-05
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100000100000100110101110100110;
		b = 32'b01001110110000101001010110100111;
		correct = 32'b00010001001010111001010110010001;
		#400 //2.2094092e-19 * 1632293800.0 = 1.353561e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100111010010010111011101001;
		b = 32'b01000111101010110010000011101000;
		correct = 32'b00111100101011100110101001011001;
		#400 //1865.466 * 87617.81 = 0.021290945
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000100010010010011101011101001;
		b = 32'b00110100110111110000010110010010;
		correct = 32'b01001110111001101111110001101100;
		#400 //804.9205 * 4.154104e-07 = 1937651200.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011101111101001010001111101100;
		b = 32'b00001101110011101010011110101000;
		correct = 32'b01001111100101111000011100011101;
		#400 //6.4755753e-21 * 1.2736092e-30 = 5084429000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00101000011111011111100101011110;
		b = 32'b10001100111111110110001001111111;
		correct = 32'b11011010111111101001011000000000;
		#400 //1.4098394e-14 * -3.934825e-31 = -3.5829785e+16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110000010011101110010100000100;
		b = 32'b00011110110001111111011011010001;
		correct = 32'b01010001000001000110111110110001;
		#400 //7.5267814e-10 * 2.1172025e-20 = 35550597000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00011010101111011100010101110110;
		b = 32'b00001111100010000100100010110011;
		correct = 32'b01001010101100100011110001110100;
		#400 //7.8487583e-23 * 1.3438638e-29 = 5840442.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110101111110000101100110011100;
		b = 32'b01100110010001101011001011001111;
		correct = 32'b10001111000111111111110000110011;
		#400 //-1.850352e-06 * 2.3458175e+23 = -7.887877e-30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100110110001110100110111101001;
		b = 32'b11100101001110011100101100100111;
		correct = 32'b00000001000010010100111011011101;
		#400 //-1.3829516e-15 * -5.483658e+22 = 2.5219508e-38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100101010000101011000100100111;
		b = 32'b10101100110010110110001000110001;
		correct = 32'b11110111111101010000111101010101;
		#400 //5.7462936e+22 * -5.7805085e-12 = -9.94081e+33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001110010001000110000001100000;
		b = 32'b10110111111110010001101101010010;
		correct = 32'b10010101110010011100111110000011;
		#400 //2.4205268e-30 * -2.9695835e-05 = -8.151065e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100001001110100000010111101110;
		b = 32'b11110011110101001110101100010110;
		correct = 32'b10101100110111111010100110110101;
		#400 //2.144701e+20 * -3.3738252e+31 = -6.3568825e-12
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000000001101100101011001101101;
		b = 32'b10101000010100111001100000011100;
		correct = 32'b11010111010111001001101010000010;
		#400 //2.849025 * -1.1745836e-14 = -242556160000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100011010010101011010111111010;
		b = 32'b00101111111011011010000010011010;
		correct = 32'b10110010110110100110001001000100;
		#400 //-1.0988977e-17 * 4.3224163e-10 = -2.5423226e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000101010011000110111001000111;
		b = 32'b01010010010000100100011000011110;
		correct = 32'b10110010100001101011000100100111;
		#400 //-3270.8923 * 208600000000.0 = -1.5680213e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010100110100101111111011111101;
		b = 32'b00111100001111011010100000010011;
		correct = 32'b11011000000011100110011011110010;
		#400 //-7249769000000.0 * 0.011575717 = -626291200000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10000101110100110111000101001111;
		b = 32'b10100100111010001100110011001001;
		correct = 32'b00100000011010001000001110100111;
		#400 //-1.9883968e-35 * -1.0096088e-16 = 1.9694724e-19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000000000100100100101010101110;
		b = 32'b00000011101110000000001010010111;
		correct = 32'b11111011110010111000011001101110;
		#400 //-2.285808 * 1.0815143e-36 = -2.1135256e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110111101001101110000011110001;
		b = 32'b01100001010111000101110010101010;
		correct = 32'b01010101110000011101110111111100;
		#400 //6.7694034e+33 * 2.5406005e+20 = 26644895000000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111011010000001010101000001100;
		b = 32'b01011110111111110111100100111011;
		correct = 32'b01011011110000010000111110101111;
		#400 //1.00036996e+36 * 9.204405e+18 = 1.0868383e+17
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110001111101011001111100100100;
		b = 32'b01001001010000110011010000101101;
		correct = 32'b00101000001000010000111101101011;
		#400 //7.1485307e-09 * 799554.8 = 8.940639e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000110000110010010001001001010;
		b = 32'b11011101110000100100111101111011;
		correct = 32'b10100111110010011100000000110011;
		#400 //9800.572 * -1.7501931e+18 = -5.599709e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100100110110011000010111011011;
		b = 32'b01110010000000111111001011000100;
		correct = 32'b00110010010100110000001110010000;
		#400 //3.210071e+22 * 2.6135054e+30 = 1.22826265e-08
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100011110110111111011111001011;
		b = 32'b00100100011110010110000111001100;
		correct = 32'b01111110111000011100111000101011;
		#400 //8.1153846e+21 * 5.4076105e-17 = 1.5007339e+38
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01011111101001000100001100111011;
		b = 32'b10111001100100001000111001110100;
		correct = 32'b11100101100100010111001011111100;
		#400 //2.3672738e+19 * -0.00027571956 = -8.585803e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111001000111101101000110101111;
		b = 32'b00101110100110110110010110101001;
		correct = 32'b11001010000000101101000110010100;
		#400 //-0.00015146167 * 7.0666424e-11 = -2143333.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111100010110010000010000010001;
		b = 32'b10011011001111101000100011101001;
		correct = 32'b01100000100100011100101000110001;
		#400 //-0.013245598 * -1.576067e-22 = 8.40421e+19
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00001010000110111011100100100111;
		b = 32'b10100001110101001100011010000101;
		correct = 32'b10100111101110110101101110011100;
		#400 //7.497802e-33 * -1.4418226e-18 = -5.200225e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10101101010010100110110100000100;
		b = 32'b01010000000000010010000011111100;
		correct = 32'b10011100110010001010011111111111;
		#400 //-1.1506577e-11 * 8665690000.0 = -1.3278316e-21
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010101010000010001001000110100;
		b = 32'b01001001110111110001001011000001;
		correct = 32'b01001010110111011001000111000011;
		#400 //13267745000000.0 * 1827416.1 = 7260385.5
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111101010100000001101000001100;
		b = 32'b00001110101110100001100111110001;
		correct = 32'b01101110000011110010000110111111;
		#400 //0.05080609 * 4.587752e-30 = 1.1074288e+28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111110001100011111101111001101;
		b = 32'b01110000101001110011100010111110;
		correct = 32'b01001101000010000011110011011101;
		#400 //5.9145195e+37 * 4.1402075e+29 = 142855630.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110101011101011110100001011110;
		b = 32'b00111000000001011110011111010011;
		correct = 32'b01111100111010110001000000000011;
		#400 //3.1172502e+32 * 3.1925574e-05 = 9.764116e+36
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01110100011101111011011100011000;
		b = 32'b10110110111000000101101001001000;
		correct = 32'b11111101000011010101010000111100;
		#400 //7.8504084e+31 * -6.6862303e-06 = -1.1741157e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010011101110110011111110001001;
		b = 32'b00101101000011010000010011100100;
		correct = 32'b01100110001010011111011000001101;
		#400 //1608449700000.0 * 8.016008e-12 = 2.006547e+23
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00111100000101010100000100111101;
		b = 32'b10110100010010000110010010111101;
		correct = 32'b11000111001111101010101111001001;
		#400 //0.009109792 * -1.86631e-07 = -48811.785
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010011001111100001101000001100;
		b = 32'b11101100010101001010000011111001;
		correct = 32'b10100110011001001110000011000010;
		#400 //816480800000.0 * -1.0282098e+27 = -7.9407994e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01001110100111010001010110001010;
		b = 32'b01111110101001110000100011011001;
		correct = 32'b00001111011100001011111111110100;
		#400 //1317717200.0 * 1.1101351e+38 = 1.18698824e-29
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110011011000000110110101010110;
		b = 32'b00000001010110101011000111000111;
		correct = 32'b11110001100000110101101011110011;
		#400 //-5.2253505e-08 * 4.0167825e-38 = -1.3008796e+30
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11011101111100001001000001000111;
		b = 32'b11010101010010110111010110111010;
		correct = 32'b01001000000101110101011110110010;
		#400 //-2.1668041e+18 * -13981656000000.0 = 154974.78
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01010000001101100111010000010111;
		b = 32'b01111000010001000010001100111110;
		correct = 32'b00010111011011100010001110101010;
		#400 //12244246000.0 * 1.5912578e+34 = 7.694696e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000110100101100010101101100101;
		b = 32'b00110101111110010001111111101001;
		correct = 32'b01010000000110100101000001011011;
		#400 //19221.697 * 1.8561233e-06 = 10355830000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010110001111100010001010001010;
		b = 32'b11101111100111111001011110101110;
		correct = 32'b00100110000110000111111100001111;
		#400 //-52263890000000.0 * -9.878297e+28 = 5.290779e-16
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11010101001011001100100111100011;
		b = 32'b11111101001111100000101101111110;
		correct = 32'b00010111011010001100000101000100;
		#400 //-11873944000000.0 * -1.5788312e+37 = 7.520718e-25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00110100111001001110111011111000;
		b = 32'b00100000010111100011001000100010;
		correct = 32'b01010100000000111110000110100000;
		#400 //4.2642182e-07 * 1.8820719e-19 = 2265704300000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001100001100111100010001101010;
		b = 32'b00100010011000001000111100111000;
		correct = 32'b11101001010011001110111110111011;
		#400 //-47124904.0 * 3.043348e-18 = -1.548456e+25
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10010010000111111111100000100101;
		b = 32'b00111100111011011011111100100100;
		correct = 32'b10010100101011000100000001001111;
		#400 //-5.0477415e-28 * 0.029021807 = -1.7392927e-26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00010111110111010011100010110100;
		b = 32'b10001111010110110000010101011111;
		correct = 32'b11001000000000010100100100111001;
		#400 //1.4296104e-24 * -1.0798568e-29 = -132388.89
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100101101110110110011110100111;
		b = 32'b00100111010110011001111010100100;
		correct = 32'b11111101110111000111010011010110;
		#400 //-1.1062432e+23 * 3.0200799e-15 = -3.66296e+37
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001101111111010000011111110000;
		b = 32'b01001101010111000110000101011001;
		correct = 32'b11000000000100101111011011001010;
		#400 //-530644480.0 * 231085460.0 = -2.2963128
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01000000111000110100101101110011;
		b = 32'b10110101011000111110111110100100;
		correct = 32'b11001010111111110100011110011000;
		#400 //7.10296 * -8.491281e-07 = -8365004.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01100011100011110001111100110110;
		b = 32'b11100010111011011011001111100010;
		correct = 32'b11000000000110100010001110001010;
		#400 //5.280267e+21 * -2.1924201e+21 = -2.4084191
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01101001001101100010010010010101;
		b = 32'b11100100011111100101011011101001;
		correct = 32'b11000100001101110101010100000010;
		#400 //1.3762328e+25 * -1.8766942e+22 = -733.32825
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100110101111011000000101110010;
		b = 32'b11011100001010000000110111001010;
		correct = 32'b10001010000100000101011011000111;
		#400 //1.3149596e-15 * -1.8921183e+17 = -6.949669e-33
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11100001011110001101000001001001;
		b = 32'b01011001100101000111000100000101;
		correct = 32'b11000111010101101000110011010111;
		#400 //-2.8686257e+20 * 5222820400000000.0 = -54924.84
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110010001100010101000100010100;
		b = 32'b01001001110010001000001001100110;
		correct = 32'b10100111111000100110001110001001;
		#400 //-1.0321191e-08 * 1642572.8 = -6.2835517e-15
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b00100111000111010001111110010011;
		b = 32'b00110001100010001111000111100101;
		correct = 32'b00110101000100101101110001000101;
		#400 //2.1805243e-15 * 3.985621e-09 = 5.470977e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b01111100100001001010101000010101;
		b = 32'b01000010100001000010110000101001;
		correct = 32'b01111001100000000111100111110010;
		#400 //5.510663e+36 * 66.08625 = 8.338592e+34
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001001111001101011010010001001;
		b = 32'b00011101111001011110011111000101;
		correct = 32'b11101011100000000111001000000001;
		#400 //-1889937.1 * 6.085544e-21 = -3.1056175e+26
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10111100100111101001101011110010;
		b = 32'b00000111011111000001101110000000;
		correct = 32'b11110100101000010000110111011100;
		#400 //-0.019360993 * 1.8966454e-34 = -1.0208019e+32
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11000000100011001011000010001010;
		b = 32'b01001011111110010001101100010101;
		correct = 32'b10110100000100001001010101010100;
		#400 //-4.39655 * 32650794.0 = -1.346537e-07
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10110001010101111011011101000010;
		b = 32'b11011110111001011010010101011010;
		correct = 32'b00010001111100000111100010101010;
		#400 //-3.1390788e-09 * -8.2738657e+18 = 3.7939688e-28
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100101000010101010100101000101;
		b = 32'b00010011101101111010000010100111;
		correct = 32'b11010000110000010100111110101110;
		#400 //-1.2026943e-16 * 4.635411e-27 = -25945797000.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b11001110010000010000111111100011;
		b = 32'b11010011101001010001001011101110;
		correct = 32'b00111010000101011011001111001000;
		#400 //-809760960.0 * -1417974400000.0 = 0.00057106884
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100010100001011010001110000000;
		b = 32'b00010110111000010101001011001100;
		correct = 32'b11001011000101111101010100110110;
		#400 //-3.6222835e-18 * 3.6402963e-25 = -9950518.0
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		a = 32'b10100110111111100010100101110111;
		b = 32'b10000001111110101110011101010000;
		correct = 32'b01100100100000011010100110001100;
		#400 //-1.763603e-15 * -9.2167413e-38 = 1.9134777e+22
					begin
			$display ("A      : %b %b %b", a[31], a[30:23], a[22:0]);
			$display ("B      : %b %b %b", b[31], b[30:23], b[22:0]);
			$display ("Output : %b %b %b", correct[31], correct[30:23], correct[22:0]);
			$display ("Correct: %b %b %b", correct[31], correct[30:23], correct[22:0]); $display();
		end

		$display ("Done.");
		$finish;
	end

endmodule